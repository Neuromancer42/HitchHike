`timescale 1 ns/100 ps
// Version: v11.8 SP2 11.8.2.4


module dbpsk_modulator(
       reset_c,
       ref_signal_c,
       whitening_0_output_whitening,
       output_data_rate_c,
       output_signal_c
    );
input  reset_c;
input  ref_signal_c;
input  whitening_0_output_whitening;
output output_data_rate_c;
input  output_signal_c;

    wire counter_n5_i_0, counter_n5_i_a3_0_0, N_123, counter_n4_i_0, 
        N_105, counter_n1_i_1, \counter[0]_net_1 , \counter_i_0[1] , 
        \counter[4]_net_1 , counter_n4_i_a3_0_0, \counter[5]_net_1 , 
        counter_n1_i_a3_0, output_dbpsk_0_sqmuxa_i_a2_8, 
        output_dbpsk_0_sqmuxa_i_a2_5, \counter[11]_net_1 , 
        \counter[12]_net_1 , output_dbpsk_0_sqmuxa_i_a2_7, 
        \counter_i_0[8] , \counter_i_0[2] , 
        output_dbpsk_0_sqmuxa_i_a2_3, output_dbpsk_0_sqmuxa_i_a2_6, 
        \counter_i_0[7] , output_dbpsk_0_sqmuxa_i_a2_1, 
        \counter[15]_net_1 , \counter[10]_net_1 , \counter[9]_net_1 , 
        \counter[14]_net_1 , \counter[13]_net_1 , \counter_i_0[6] , 
        \counter_i_0[3] , output_dbpsk_0_sqmuxa_i_a3_2, 
        output_dbpsk_0_sqmuxa_i_a3_1, N_122, 
        output_dbpsk_0_sqmuxa_i_a3_0, N_11, N_35, N_13, N_34, N_15, 
        N_33, N_21, N_30, N_23, N_29, N_25, N_19, N_32, N_106, N_17, 
        output_dbpsk_5, counter_n0, counter_n15, N_42, counter_n14, 
        N_41, counter_n13, N_40, counter_n12, N_39, counter_n11, N_38, 
        counter_n10, N_37, counter_n9, N_36, N_28, GND, VCC;
    
    NOR3B \counter_RNI29ND[15]  (.A(\counter_i_0[7] ), .B(
        output_dbpsk_0_sqmuxa_i_a2_1), .C(\counter[15]_net_1 ), .Y(
        output_dbpsk_0_sqmuxa_i_a2_6));
    NOR2 output_dbpsk_RNO_3 (.A(\counter[4]_net_1 ), .B(
        \counter[5]_net_1 ), .Y(output_dbpsk_0_sqmuxa_i_a3_0));
    XAI1A \counter_RNO_1[1]  (.A(\counter[0]_net_1 ), .B(
        \counter_i_0[1] ), .C(output_signal_c), .Y(counter_n1_i_1));
    XA1A \counter_RNO[12]  (.A(\counter[12]_net_1 ), .B(N_39), .C(
        output_signal_c), .Y(counter_n12));
    DFN1E1C0 output_dbpsk (.D(output_dbpsk_5), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(N_28), .Q(output_data_rate_c));
    DFN1P0 \counter[2]  (.D(N_23), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\counter_i_0[2] ));
    NOR3B output_dbpsk_RNO_2 (.A(\counter_i_0[1] ), .B(
        output_dbpsk_0_sqmuxa_i_a3_0), .C(\counter[0]_net_1 ), .Y(
        output_dbpsk_0_sqmuxa_i_a3_1));
    DFN1P0 \counter[7]  (.D(N_13), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\counter_i_0[7] ));
    NOR2B \counter_RNO_2[4]  (.A(\counter_i_0[1] ), .B(
        \counter[5]_net_1 ), .Y(counter_n4_i_a3_0_0));
    NOR2A \counter_RNO[0]  (.A(output_signal_c), .B(\counter[0]_net_1 )
        , .Y(counter_n0));
    DFN1P0 \counter[6]  (.D(N_15), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\counter_i_0[6] ));
    NOR3A \counter_RNO[4]  (.A(N_32), .B(N_106), .C(counter_n4_i_0), 
        .Y(N_19));
    VCC VCC_i (.Y(VCC));
    OR2 \counter_RNIGL45[2]  (.A(\counter_i_0[2] ), .B(N_29), .Y(N_30));
    DFN1P0 \counter[8]  (.D(N_11), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\counter_i_0[8] ));
    AO1B output_dbpsk_RNO_0 (.A(output_dbpsk_0_sqmuxa_i_a3_2), .B(
        whitening_0_output_whitening), .C(output_signal_c), .Y(N_28));
    NOR2B \counter_RNO_0[1]  (.A(\counter[4]_net_1 ), .B(
        \counter[5]_net_1 ), .Y(counter_n1_i_a3_0));
    AO1 \counter_RNO[1]  (.A(counter_n1_i_a3_0), .B(N_123), .C(
        counter_n1_i_1), .Y(N_25));
    DFN1C0 \counter[15]  (.D(counter_n15), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[15]_net_1 ));
    OR2A \counter_RNI32OP[10]  (.A(\counter[10]_net_1 ), .B(N_37), .Y(
        N_38));
    OR2A \counter_RNI316H[9]  (.A(\counter[9]_net_1 ), .B(N_36), .Y(
        N_37));
    DFN1C0 \counter[14]  (.D(counter_n14), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[14]_net_1 ));
    NOR2B \counter_RNI70E3[6]  (.A(\counter_i_0[6] ), .B(
        \counter_i_0[3] ), .Y(output_dbpsk_0_sqmuxa_i_a2_1));
    XAI1 \counter_RNO[8]  (.A(N_35), .B(\counter_i_0[8] ), .C(
        output_signal_c), .Y(N_11));
    XA1A \counter_RNO[14]  (.A(\counter[14]_net_1 ), .B(N_41), .C(
        output_signal_c), .Y(counter_n14));
    XA1A \counter_RNO[11]  (.A(\counter[11]_net_1 ), .B(N_38), .C(
        output_signal_c), .Y(counter_n11));
    DFN1C0 \counter[4]  (.D(N_19), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[4]_net_1 ));
    OA1B \counter_RNO_3[4]  (.A(N_30), .B(\counter_i_0[3] ), .C(
        \counter[4]_net_1 ), .Y(N_105));
    OR2A \counter_RNIVND3[0]  (.A(\counter[0]_net_1 ), .B(
        \counter_i_0[1] ), .Y(N_29));
    DFN1C0 \counter[5]  (.D(N_17), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[5]_net_1 ));
    OR2A \counter_RNI9BEJ1[13]  (.A(\counter[13]_net_1 ), .B(N_40), .Y(
        N_41));
    NOR2 \counter_RNI794H[13]  (.A(\counter[14]_net_1 ), .B(
        \counter[13]_net_1 ), .Y(output_dbpsk_0_sqmuxa_i_a2_3));
    XAI1 \counter_RNO[2]  (.A(N_29), .B(\counter_i_0[2] ), .C(
        output_signal_c), .Y(N_23));
    NOR2B \counter_RNO_1[5]  (.A(\counter_i_0[1] ), .B(
        \counter[4]_net_1 ), .Y(counter_n5_i_a3_0_0));
    GND GND_i (.Y(GND));
    XA1C \counter_RNO[5]  (.A(\counter[5]_net_1 ), .B(N_32), .C(
        counter_n5_i_0), .Y(N_17));
    XAI1 \counter_RNO[3]  (.A(N_30), .B(\counter_i_0[3] ), .C(
        output_signal_c), .Y(N_21));
    DFN1C0 \counter[12]  (.D(counter_n12), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[12]_net_1 ));
    DFN1P0 \counter[1]  (.D(N_25), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\counter_i_0[1] ));
    OR2 \counter_RNIKOND[7]  (.A(\counter_i_0[7] ), .B(N_34), .Y(N_35));
    AO1B \counter_RNO_0[5]  (.A(counter_n5_i_a3_0_0), .B(N_123), .C(
        output_signal_c), .Y(counter_n5_i_0));
    OR2 \counter_RNIUL0C[6]  (.A(\counter_i_0[6] ), .B(N_33), .Y(N_34));
    DFN1P0 \counter[3]  (.D(N_21), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\counter_i_0[3] ));
    XAI1 \counter_RNO[6]  (.A(N_33), .B(\counter_i_0[6] ), .C(
        output_signal_c), .Y(N_15));
    NOR3A \counter_RNIRADR[11]  (.A(output_dbpsk_0_sqmuxa_i_a2_5), .B(
        \counter[11]_net_1 ), .C(\counter[12]_net_1 ), .Y(
        output_dbpsk_0_sqmuxa_i_a2_8));
    OR3A \counter_RNILJI8[3]  (.A(\counter[4]_net_1 ), .B(N_30), .C(
        \counter_i_0[3] ), .Y(N_32));
    NOR2B output_dbpsk_RNO_1 (.A(output_dbpsk_0_sqmuxa_i_a3_1), .B(
        N_122), .Y(output_dbpsk_0_sqmuxa_i_a3_2));
    XA1A \counter_RNO[13]  (.A(\counter[13]_net_1 ), .B(N_40), .C(
        output_signal_c), .Y(counter_n13));
    OR2 \counter_RNIBSEF[8]  (.A(\counter_i_0[8] ), .B(N_35), .Y(N_36));
    XA1A \counter_RNO[9]  (.A(\counter[9]_net_1 ), .B(N_36), .C(
        output_signal_c), .Y(counter_n9));
    OR2A \counter_RNI44A21[11]  (.A(\counter[11]_net_1 ), .B(N_38), .Y(
        N_39));
    OR2A \counter_RNI9K9A[5]  (.A(\counter[5]_net_1 ), .B(N_32), .Y(
        N_33));
    NOR3C \counter_RNICUMT1[2]  (.A(output_dbpsk_0_sqmuxa_i_a2_7), .B(
        output_dbpsk_0_sqmuxa_i_a2_6), .C(output_dbpsk_0_sqmuxa_i_a2_8)
        , .Y(N_122));
    DFN1C0 \counter[11]  (.D(counter_n11), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[11]_net_1 ));
    OR2A \counter_RNO_0[15]  (.A(\counter[14]_net_1 ), .B(N_41), .Y(
        N_42));
    XA1A \counter_RNO[15]  (.A(\counter[15]_net_1 ), .B(N_42), .C(
        output_signal_c), .Y(counter_n15));
    OR2A \counter_RNO_1[4]  (.A(output_signal_c), .B(N_105), .Y(
        counter_n4_i_0));
    NOR2B \counter_RNO_0[4]  (.A(counter_n4_i_a3_0_0), .B(N_123), .Y(
        N_106));
    NOR2B \counter_RNIRPDV1[0]  (.A(N_122), .B(\counter[0]_net_1 ), .Y(
        N_123));
    OR2A \counter_RNI67SA1[12]  (.A(\counter[12]_net_1 ), .B(N_39), .Y(
        N_40));
    XAI1 \counter_RNO[7]  (.A(N_34), .B(\counter_i_0[7] ), .C(
        output_signal_c), .Y(N_13));
    NOR2A output_dbpsk_RNO (.A(output_signal_c), .B(output_data_rate_c)
        , .Y(output_dbpsk_5));
    XA1A \counter_RNO[10]  (.A(\counter[10]_net_1 ), .B(N_37), .C(
        output_signal_c), .Y(counter_n10));
    DFN1C0 \counter[13]  (.D(counter_n13), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[13]_net_1 ));
    NOR2 \counter_RNIO59A[9]  (.A(\counter[10]_net_1 ), .B(
        \counter[9]_net_1 ), .Y(output_dbpsk_0_sqmuxa_i_a2_5));
    NOR3C \counter_RNIFAIK[2]  (.A(\counter_i_0[8] ), .B(
        \counter_i_0[2] ), .C(output_dbpsk_0_sqmuxa_i_a2_3), .Y(
        output_dbpsk_0_sqmuxa_i_a2_7));
    DFN1C0 \counter[0]  (.D(counter_n0), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[0]_net_1 ));
    DFN1C0 \counter[10]  (.D(counter_n10), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[10]_net_1 ));
    DFN1C0 \counter[9]  (.D(counter_n9), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[9]_net_1 ));
    
endmodule


module randgen(
       randgen_0_cur_rand,
       ref_signal_c,
       reset_c
    );
output [23:3] randgen_0_cur_rand;
input  ref_signal_c;
input  reset_c;

    wire \mult1_un26_sum[4] , I2_un1_CO1, I3_un3_CO1, N85, 
        \rd[22]_net_1 , \rd[21]_net_1 , \mult1_un26_sum[2] , 
        \mult1_un19_sum[1] , ADD_5x5_slow_I4_Y_1, I2_un1_CO1_0, 
        \mult1_un19_sum[2] , \DWACT_ADD_CI_0_g_array_1[0] , 
        \DWACT_ADD_CI_0_TMP[0] , ADD_5x5_slow_I1_S, N85_0, 
        \rd[23]_net_1 , ADD_5x5_slow_I2_un1_CO1_0, I1_un3_CO1, 
        \mult1_un19_sum_0[1] , N74, \mult1_un19_sum_0[2] , N85_1, 
        \mult1_un19_sum_1[1] , ADD_5x5_slow_I4_Y_2, 
        ADD_5x5_slow_I4_Y_1_0, \mult1_un75_sum[4] , 
        \mult1_un89_sum[4] , N89, ADD_5x5_slow_I4_Y_2_0, N85_2, 
        I1_un2_CO1, ADD_5x5_slow_I1_CO1_0, \mult1_un82_sum[4] , N89_0, 
        I2_un1_CO1_1, I2_un1_CO1_1_tz, \mult1_un145_sum[1] , 
        \mult1_un145_sum[4] , I3_un3_CO1_0, ADD_5x5_slow_I3_CO1_0, 
        I3_un3_CO1_1, ADD_5x5_slow_I3_CO1_0_0, ADD_5x5_slow_I4_Y_1_1, 
        \mult1_un82_sum_0[4] , ADD_5x5_slow_I4_Y_2_1, I2_un1_CO1_2, 
        ADD_5x5_slow_I4_Y_0, \mult1_un166_sum[4] , 
        \mult1_un159_sum[2] , \mult1_un159_sum[4] , 
        ADD_5x5_slow_I2_S_0, ADD_4x4_slow_I1_S_0, 
        ADD_5x5_slow_I1_CO1_0_0, \rd[1]_net_1 , \rd[0]_net_1 , 
        ADD_5x5_slow_I4_Y_2_2, I2_un1_CO1_3, ADD_5x5_slow_I4_Y_0_0, 
        \mult1_un152_sum[2] , \mult1_un152_sum[4] , 
        ADD_5x5_slow_I2_S_0_0, \mult1_un159_sum[1] , 
        ADD_5x5_slow_I1_CO1_0_1, \rd[2]_net_1 , ADD_5x5_slow_I4_Y_2_3, 
        I2_un1_CO1_4, ADD_5x5_slow_I4_Y_0_1, \mult1_un166_sum_0[4] , 
        \mult1_un159_sum_0[2] , \mult1_un159_sum_0[4] , 
        ADD_5x5_slow_I4_Y_2_4, I2_un1_CO1_5, ADD_5x5_slow_I4_Y_0_2, 
        \mult1_un145_sum[2] , \mult1_un145_sum_0[4] , 
        ADD_5x5_slow_I2_S_0_1, \mult1_un166_sum[1] , 
        ADD_5x5_slow_I1_CO1_0_2, ADD_5x5_slow_I2_S_0_2, 
        \mult1_un152_sum[1] , ADD_5x5_slow_I4_Y_2_5, I2_un1_CO1_6, 
        ADD_5x5_slow_I4_Y_0_3, \mult1_un152_sum_0[2] , 
        \mult1_un152_sum_0[4] , ADD_5x5_slow_I1_CO1_0_3, \rd[3]_net_1 , 
        ADD_5x5_slow_I4_Y_2_6, I2_un1_CO1_7, ADD_5x5_slow_I4_Y_0_4, 
        \mult1_un138_sum[2] , \mult1_un138_sum[4] , 
        ADD_5x5_slow_I4_Y_2_7, I2_un1_CO1_8, ADD_5x5_slow_I4_Y_0_5, 
        \mult1_un145_sum_0[2] , ADD_5x5_slow_I4_Y_2_8, I2_un1_CO1_9, 
        ADD_5x5_slow_I4_Y_0_6, \mult1_un131_sum[2] , 
        \mult1_un131_sum[4] , ADD_5x5_slow_I2_S_0_3, 
        \mult1_un138_sum[1] , ADD_5x5_slow_I4_Y_2_9, I2_un1_CO1_10, 
        ADD_5x5_slow_I4_Y_0_7, \mult1_un138_sum_0[2] , 
        \mult1_un138_sum_0[4] , ADD_5x5_slow_I4_Y_2_10, I2_un1_CO1_11, 
        ADD_5x5_slow_I4_Y_0_8, \mult1_un124_sum[2] , 
        \mult1_un124_sum[4] , ADD_5x5_slow_I2_S_0_4, \rd[4]_net_1 , 
        ADD_5x5_slow_I4_Y_2_11, I2_un1_CO1_12, ADD_5x5_slow_I4_Y_0_9, 
        \mult1_un131_sum_0[2] , \mult1_un131_sum_0[4] , 
        ADD_5x5_slow_I4_Y_2_12, I2_un1_CO1_13, ADD_5x5_slow_I4_Y_0_10, 
        \mult1_un117_sum[2] , \mult1_un117_sum[4] , 
        ADD_5x5_slow_I2_S_0_5, \mult1_un138_sum_0[1] , 
        ADD_5x5_slow_I4_Y_2_13, I2_un1_CO1_14, ADD_5x5_slow_I4_Y_0_11, 
        \mult1_un124_sum_0[2] , \mult1_un124_sum_0[4] , 
        ADD_5x5_slow_I4_Y_2_14, I2_un1_CO1_15, ADD_5x5_slow_I4_Y_0_12, 
        \mult1_un110_sum[2] , \mult1_un110_sum[4] , 
        ADD_5x5_slow_I4_Y_2_15, I2_un1_CO1_16, ADD_5x5_slow_I4_Y_0_13, 
        \mult1_un117_sum_0[2] , \mult1_un117_sum_0[4] , 
        ADD_4x4_slow_I3_Y_1, I1_un2_CO1_0, ADD_4x4_slow_I1_CO1_0, 
        ADD_4x4_slow_I3_Y_0, \mult1_un159_sum_0[1] , 
        \mult1_un159_sum[3] , ADD_5x5_slow_I4_Y_2_16, 
        ADD_5x5_slow_I4_Y_1_2, \mult1_un103_sum[4] , 
        \mult1_un103_sum[2] , I2_un1_CO1_17, ADD_4x4_slow_I3_Y_2, 
        N74_0, ADD_4x4_slow_I3_Y_0_0, I2_un1_CO1_18, 
        ADD_4x4_slow_I3_Y_2_0, \mult1_un152_sum_0[1] , 
        ADD_5x5_slow_I4_Y_2_17, ADD_5x5_slow_I4_Y_1_3, I2_un1_CO1_1_0, 
        I2_un5_CO1, ADD_5x5_slow_I4_Y_0_14, \mult1_un110_sum_0[2] , 
        \mult1_un110_sum_0[4] , ADD_5x5_slow_I2_S_0_6, 
        \mult1_un110_sum[1] , ADD_4x4_slow_I3_Y_2_1, 
        ADD_4x4_slow_I3_Y_1_0, ADD_4x4_slow_I3_Y_0_1, N74_1, 
        \mult1_un138_sum[3] , ADD_4x4_slow_I1_S_0_0, 
        \mult1_un145_sum[3] , ADD_5x5_slow_I4_Y_2_18, 
        ADD_5x5_slow_I4_Y_1_4, \mult1_un96_sum[4] , 
        \mult1_un96_sum[2] , I2_un1_CO1_19, ADD_5x5_slow_I4_Y_2_19, 
        I2_un1_CO1_20, ADD_5x5_slow_I4_Y_0_15, \mult1_un103_sum_0[2] , 
        \mult1_un103_sum_0[4] , ADD_4x4_slow_I1_S_0_1, 
        ADD_5x5_slow_I2_S_0_7, \mult1_un103_sum[1] , N74_2, 
        ADD_4x4_slow_I3_Y_0_2, \mult1_un138_sum_1[1] , 
        ADD_5x5_slow_I4_Y_2_20, I2_un1_CO1_21, ADD_5x5_slow_I4_Y_0_16, 
        \mult1_un89_sum[2] , ADD_4x4_slow_I1_CO1_0_0, 
        ADD_4x4_slow_I1_S_0_2, ADD_5x5_slow_I4_Y_2_21, 
        ADD_5x5_slow_I4_Y_1_5, \mult1_un96_sum_0[4] , 
        \mult1_un96_sum_0[2] , I2_un1_CO1_22, ADD_4x4_slow_I3_Y_2_2, 
        N74_3, ADD_4x4_slow_I3_Y_0_3, \mult1_un131_sum[1] , 
        \mult1_un131_sum[3] , ADD_4x4_slow_I1_CO1_0_1, \rd[5]_net_1 , 
        ADD_4x4_slow_I3_Y_2_3, ADD_4x4_slow_I3_Y_1_1, 
        ADD_4x4_slow_I3_Y_0_4, N74_4, \mult1_un124_sum[1] , 
        \mult1_un124_sum[3] , ADD_5x5_slow_I4_Y_2_22, I2_un1_CO1_23, 
        ADD_5x5_slow_I4_Y_0_17, \mult1_un82_sum[2] , 
        ADD_5x5_slow_I4_Y_2_23, I2_un1_CO1_24, ADD_5x5_slow_I4_Y_0_18, 
        \mult1_un89_sum_0[2] , \mult1_un89_sum_0[4] , 
        ADD_4x4_slow_I1_S_0_3, \rd[6]_net_1 , ADD_4x4_slow_I3_Y_2_4, 
        ADD_4x4_slow_I3_Y_1_2, \mult1_un117_sum[3] , 
        \mult1_un117_sum[1] , N74_5, ADD_5x5_slow_I4_Y_2_24, 
        I2_un1_CO1_25, ADD_5x5_slow_I4_Y_0_19, \mult1_un82_sum_0[2] , 
        \mult1_un75_sum_0[4] , \mult1_un75_sum[2] , I2_un1_CO1_26, 
        ADD_4x4_slow_I1_S_0_4, \rd[7]_net_1 , ADD_4x4_slow_I3_Y_2_5, 
        ADD_4x4_slow_I3_Y_1_3, \mult1_un110_sum[3] , 
        \mult1_un110_sum_0[1] , N74_6, ADD_5x5_slow_I2_S_0_8, 
        \mult1_un82_sum[1] , ADD_5x5_slow_I4_Y_2_25, I2_un1_CO1_27, 
        ADD_5x5_slow_I4_Y_0_20, \mult1_un75_sum_0[2] , 
        ADD_4x4_slow_I1_S_0_5, \rd[8]_net_1 , ADD_4x4_slow_I3_Y_2_6, 
        ADD_4x4_slow_I3_Y_1_4, \mult1_un103_sum[3] , 
        \mult1_un103_sum_0[1] , N74_7, ADD_5x5_slow_I4_Y_2_26, 
        I2_un1_CO1_28, ADD_5x5_slow_I4_Y_0_21, \mult1_un68_sum[2] , 
        \mult1_un68_sum[4] , ADD_5x5_slow_I2_S_0_9, 
        \mult1_un75_sum[1] , ADD_4x4_slow_I1_S_0_6, \rd[9]_net_1 , 
        I2_un1_CO1_1_1, I2_un5_CO1_0, ADD_5x5_slow_I4_Y_0_22, 
        \mult1_un68_sum_0[2] , \mult1_un68_sum_0[4] , 
        ADD_5x5_slow_I1_CO1_0_4, \rd[14]_net_1 , \rd[13]_net_1 , 
        ADD_4x4_slow_I3_Y_2_7, ADD_4x4_slow_I3_Y_1_5, 
        \mult1_un96_sum[3] , \mult1_un96_sum[1] , N74_8, 
        ADD_5x5_slow_I4_Y_2_27, I2_un1_CO1_29, ADD_5x5_slow_I4_Y_0_23, 
        \mult1_un61_sum[2] , \mult1_un61_sum[4] , 
        ADD_5x5_slow_I2_S_0_10, \mult1_un75_sum_0[1] , 
        ADD_4x4_slow_I1_S_0_7, \rd[10]_net_1 , ADD_5x5_slow_I1_CO1_0_5, 
        ADD_4x4_slow_I3_Y_2_8, ADD_4x4_slow_I3_Y_1_6, 
        \mult1_un89_sum[3] , \mult1_un89_sum[1] , N74_9, 
        ADD_5x5_slow_I2_S_2, N83, ADD_5x5_slow_I2_S_2_0, 
        ADD_5x5_slow_I2_S_1, \mult1_un152_sum[3] , 
        ADD_5x5_slow_I4_Y_2_28, ADD_5x5_slow_I4_Y_1_6, 
        \mult1_un61_sum_0[4] , \mult1_un61_sum_0[2] , I2_un1_CO1_30, 
        ADD_4x4_slow_I1_S_0_8, \rd[11]_net_1 , ADD_5x5_slow_I2_S_1_0, 
        \mult1_un145_sum_0[3] , ADD_5x5_slow_I4_Y_2_29, 
        ADD_5x5_slow_I4_Y_1_7, \mult1_un54_sum[4] , 
        \mult1_un54_sum[2] , I2_un1_CO1_31, ADD_4x4_slow_I3_Y_2_9, 
        N74_10, ADD_4x4_slow_I3_Y_0_5, \mult1_un82_sum_0[1] , 
        \mult1_un82_sum[3] , ADD_5x5_slow_I2_S_2_1, 
        ADD_5x5_slow_I2_S_1_1, \mult1_un138_sum_0[3] , 
        ADD_5x5_slow_I4_Y_2_30, ADD_5x5_slow_I4_Y_1_8, I2_un1_CO1_1_2, 
        I2_un5_CO1_1, ADD_5x5_slow_I4_Y_0_24, \mult1_un54_sum_0[2] , 
        \mult1_un54_sum_0[4] , ADD_4x4_slow_I1_S_0_9, \rd[12]_net_1 , 
        ADD_4x4_slow_I3_Y_2_10, N74_11, ADD_4x4_slow_I3_Y_0_6, 
        \mult1_un75_sum_1[1] , \mult1_un75_sum[3] , 
        ADD_5x5_slow_I2_S_2_2, ADD_5x5_slow_I2_S_1_2, 
        \mult1_un131_sum_0[3] , ADD_5x5_slow_I4_Y_2_31, 
        ADD_5x5_slow_I4_Y_1_9, \mult1_un47_sum[4] , 
        \mult1_un47_sum[2] , I2_un1_CO1_32, ADD_4x4_slow_I1_S_0_10, 
        ADD_5x5_slow_I2_S_2_3, ADD_5x5_slow_I2_S_1_3, 
        \mult1_un124_sum_0[3] , ADD_4x4_slow_I3_Y_2_11, N74_12, 
        ADD_4x4_slow_I3_Y_0_7, \mult1_un68_sum[1] , 
        \mult1_un68_sum[3] , ADD_5x5_slow_I4_Y_2_32, I2_un1_CO1_33, 
        ADD_5x5_slow_I4_Y_0_25, \mult1_un47_sum_0[2] , 
        \mult1_un47_sum_0[4] , ADD_5x5_slow_I2_S_2_4, 
        ADD_5x5_slow_I2_S_1_4, \mult1_un117_sum_0[3] , 
        ADD_4x4_slow_I1_CO1_0_2, ADD_4x4_slow_I1_S_0_11, 
        ADD_5x5_slow_I4_Y_2_33, ADD_5x5_slow_I4_Y_1_10, 
        \mult1_un40_sum[4] , \mult1_un40_sum[2] , I2_un1_CO1_34, 
        ADD_4x4_slow_I3_Y_2_12, ADD_4x4_slow_I3_Y_1_7, 
        \mult1_un61_sum[3] , \mult1_un61_sum[1] , N74_13, 
        ADD_5x5_slow_I2_S_2_5, ADD_5x5_slow_I2_S_1_5, 
        \mult1_un110_sum_0[3] , ADD_5x5_slow_I4_Y_2_34, 
        ADD_5x5_slow_I4_Y_1_11, \mult1_un40_sum_0[4] , 
        \mult1_un40_sum_0[2] , I2_un1_CO1_35, ADD_4x4_slow_I1_S_0_12, 
        \rd[15]_net_1 , ADD_5x5_slow_I2_S_2_6, ADD_5x5_slow_I2_S_1_6, 
        \mult1_un103_sum_0[3] , ADD_4x4_slow_I3_Y_2_13, N74_14, 
        ADD_4x4_slow_I3_Y_0_8, \mult1_un54_sum[1] , 
        \mult1_un54_sum[3] , ADD_5x5_slow_I2_S_2_7, 
        ADD_5x5_slow_I2_S_1_7, \mult1_un96_sum_0[3] , 
        ADD_5x5_slow_I4_Y_2_35, ADD_5x5_slow_I4_Y_1_12, 
        \mult1_un33_sum[4] , \mult1_un33_sum[2] , I2_un1_CO1_36, 
        ADD_4x4_slow_I1_S_0_13, \rd[16]_net_1 , ADD_5x5_slow_I4_Y_2_36, 
        ADD_5x5_slow_I4_Y_1_13, \mult1_un33_sum_0[4] , 
        \mult1_un33_sum_0[2] , I2_un1_CO1_37, ADD_4x4_slow_I3_Y_2_14, 
        N74_15, ADD_4x4_slow_I3_Y_0_9, \mult1_un47_sum[1] , 
        \mult1_un47_sum[3] , ADD_5x5_slow_I2_S_2_8, 
        ADD_5x5_slow_I2_S_1_8, \mult1_un89_sum_0[3] , 
        ADD_5x5_slow_I2_S_2_9, ADD_5x5_slow_I2_S_1_9, N83_0, 
        ADD_5x5_slow_I2_S_2_10, ADD_4x4_slow_I1_S_0_14, \rd[17]_net_1 , 
        ADD_5x5_slow_I4_Y_2_37, I2_un1_CO1_38, ADD_5x5_slow_I4_Y_0_26, 
        ADD_4x4_slow_I3_Y_2_15, N74_16, ADD_4x4_slow_I3_Y_0_10, 
        \mult1_un40_sum[1] , \mult1_un40_sum[3] , 
        ADD_5x5_slow_I4_Y_2_38, ADD_5x5_slow_I4_Y_1_14, 
        \mult1_un26_sum_0[4] , \mult1_un26_sum_0[2] , I2_un1_CO1_39, 
        ADD_5x5_slow_I2_S_2_11, ADD_5x5_slow_I2_S_1_10, 
        \mult1_un75_sum_0[3] , ADD_4x4_slow_I1_S_0_15, \rd[18]_net_1 , 
        ADD_5x5_slow_I2_S_1_11, \mult1_un68_sum_0[3] , 
        ADD_4x4_slow_I3_Y_2_16, ADD_4x4_slow_I3_Y_1_8, 
        \mult1_un33_sum[3] , \mult1_un33_sum[1] , N74_17, 
        ADD_5x5_slow_I4_Y_2_39, ADD_5x5_slow_I2_S_2_12, 
        ADD_5x5_slow_I2_S_1_12, \mult1_un61_sum_0[3] , 
        ADD_5x5_slow_I4_Y_2_40, ADD_5x5_slow_I4_Y_1_15, 
        \mult1_un19_sum[4] , I2_un1_CO1_40, ADD_4x4_slow_I1_S_0_16, 
        \rd[19]_net_1 , ADD_4x4_slow_I3_Y_2_17, ADD_4x4_slow_I3_Y_1_9, 
        \mult1_un26_sum[3] , \mult1_un26_sum[1] , N74_18, 
        ADD_5x5_slow_I2_S_2_13, ADD_5x5_slow_I2_S_1_13, 
        \mult1_un54_sum_0[3] , ADD_4x4_slow_I1_S_0_17, \rd[20]_net_1 , 
        ADD_5x5_slow_I2_S_2_14, ADD_5x5_slow_I2_S_1_14, 
        \mult1_un47_sum_0[3] , ADD_5x5_slow_I4_Y_2_41, 
        ADD_5x5_slow_I4_Y_1_16, I2_un4_CO1, ADD_4x4_slow_I3_Y_2_18, 
        ADD_4x4_slow_I3_Y_1_10, \mult1_un19_sum[3] , N74_19, 
        ADD_5x5_slow_I2_S_2_15, ADD_5x5_slow_I2_S_1_15, 
        \mult1_un40_sum_1[4] , ADD_4x4_slow_I1_S_0_18, 
        ADD_4x4_slow_I3_Y_2_19, ADD_5x5_slow_I2_S_2_16, 
        ADD_5x5_slow_I2_S_1_16, I2_un4_CO1_0, ADD_4x4_slow_I1_S_0_19, 
        ADD_5x5_slow_I2_S_3, N89_1, N85_3, N85_4, I3_un3_CO1_2, 
        ADD_5x5_slow_I3_CO1_0_1, N85_5, I3_un3_CO1_3, 
        ADD_5x5_slow_I3_CO1_0_2, \mult1_un61_sum_0[1] , N85_6, 
        I3_un3_CO1_4, ADD_5x5_slow_I3_CO1_0_3, \mult1_un68_sum_0[1] , 
        N85_7, I1_un2_CO1_1, I1_un5_CO1, I1_un3_CO1_0, I1_un2_CO1_2, 
        \mult1_un89_sum_0[1] , N85_8, N85_9, \mult1_un96_sum_0[1] , 
        N85_10, N85_11, \mult1_un47_sum_0[1] , N83_1, 
        \mult1_un33_sum_0[1] , I2_un4_CO1_1, ADD_4x4_slow_I2_un1_CO1_0, 
        I2_un4_CO1_2, ADD_4x4_slow_I2_un1_CO1_0_0, I1_un2_CO1_3, 
        N85_12, N85_13, N89_2, N89_3, I3_un3_CO1_5, 
        ADD_5x5_slow_I3_CO1_0_4, N85_14, I3_un3_CO1_6, 
        ADD_5x5_slow_I3_CO1_0_5, \mult1_un40_sum_0[1] , 
        \mult1_un54_sum_0[1] , I2_un4_CO1_3, 
        ADD_4x4_slow_I2_un1_CO1_0_1, N89_4, N83_2, N83_3, I3_un3_CO1_7, 
        ADD_5x5_slow_I3_CO1_0_6, \mult1_un131_sum_0[1] , N85_15, 
        \mult1_un124_sum_0[1] , N83_4, I3_un3_CO1_8, 
        ADD_5x5_slow_I3_CO1_0_7, \mult1_un131_sum_1[1] , N85_16, 
        I3_un3_CO1_9, ADD_5x5_slow_I3_CO1_0_8, I3_un3_CO1_10, 
        ADD_5x5_slow_I3_CO1_0_9, \mult1_un117_sum_0[1] , N85_17, 
        I2_un4_CO1_4, ADD_4x4_slow_I2_un1_CO1_0_2, I2_un4_CO1_5, 
        ADD_4x4_slow_I2_un1_CO1_0_3, I1_un2_CO1_4, I1_un2_CO1_5, 
        I3_un3_CO1_11, ADD_5x5_slow_I3_CO1_0_10, I3_un3_CO1_12, 
        ADD_5x5_slow_I3_CO1_0_11, \mult1_un166_sum[2] , N85_18, 
        ADD_5x5_slow_I4_Y_0_27, I3_un3_CO1_13, 
        ADD_5x5_slow_I3_CO1_0_12, I1_un2_CO1_6, ADD_5x5_slow_I2_S_0_11, 
        I1_un2_CO1_7, ADD_5x5_slow_I1_S_1, N85_19, I3_un3_CO1_14, 
        ADD_5x5_slow_I3_CO1_0_13, ADD_5x5_slow_I4_Y, I3_un3_CO1_15, 
        ADD_5x5_slow_I3_CO1_0_14, N85_20, I2_un4_CO1_6, 
        ADD_4x4_slow_I2_un1_CO1_0_4, \mult1_un166_sum[3] , 
        I2_un4_CO1_7, ADD_4x4_slow_I2_un1_CO1_0_5, ADD_4x4_slow_I3_Y, 
        I2_un1_CO1_41, N74_20, ADD_4x4_slow_I1_S, 
        \mult1_un166_sum_0[1] , I3_un3_CO1_16, 
        ADD_5x5_slow_I3_CO1_0_15, N85_21, I1_un2_CO1_8, 
        \mult1_un145_sum_0[1] , \mult1_un124_sum_1[1] , N85_22, 
        I3_un3_CO1_17, ADD_5x5_slow_I3_CO1_0_16, I3_un3_CO1_18, 
        ADD_5x5_slow_I3_CO1_0_17, N85_23, I3_un3_CO1_19, 
        ADD_5x5_slow_I3_CO1_0_18, \mult1_un117_sum_1[1] , N85_24, 
        N89_5, I2_un1_CO1_42, N89_6, N83_5, N85_25, N85_26, N83_6, 
        I3_un3_CO1_20, ADD_5x5_slow_I3_CO1_0_19, 
        \mult1_un110_sum_1[1] , N85_27, N83_7, I3_un3_CO1_21, 
        ADD_5x5_slow_I3_CO1_0_20, N83_8, N83_9, N83_10, N83_11, 
        I2_un1_CO1_43, I2_un4_CO1_8, ADD_4x4_slow_I2_un1_CO1_0_6, 
        N85_28, N83_12, I1_un5_CO1_0, I1_un3_CO1_1, I1_un2_CO1_9, 
        I3_un3_CO1_22, ADD_5x5_slow_I3_CO1_0_21, \mult1_un54_sum_1[1] , 
        N85_29, N89_7, \mult1_un68_sum_1[1] , N85_30, N89_8, 
        I3_un3_CO1_23, ADD_5x5_slow_I3_CO1_0_22, \mult1_un40_sum_1[1] , 
        \mult1_un47_sum_1[1] , N85_31, I1_un2_CO1_10, 
        \mult1_un82_sum_1[1] , I3_un3_CO1_24, ADD_5x5_slow_I3_CO1_0_23, 
        \mult1_un61_sum_1[1] , N85_32, I3_un3_CO1_25, 
        ADD_5x5_slow_I3_CO1_0_24, I3_un3_CO1_26, 
        ADD_5x5_slow_I3_CO1_0_25, \mult1_un26_sum_0[1] , N85_33, 
        \mult1_un33_sum_1[1] , N85_34, I3_un3_CO1_27, 
        ADD_5x5_slow_I3_CO1_0_26, N83_13, N83_14, I1_un5_CO1_1, 
        I1_un3_CO1_2, I1_un2_CO1_11, ADD_5x5_slow_I1_S_0, N83_15, 
        I1_un5_CO1_2, I1_un3_CO1_3, I1_un2_CO1_12, 
        \mult1_un166_sum_0[2] , \mult1_un166_sum_1[2] , 
        \mult1_un159_sum_1[1] , ADD_5x5_slow_I2_S, N85_35, 
        I3_un3_CO1_28, ADD_5x5_slow_I3_CO1_0_27, 
        \mult1_un152_sum_1[1] , N85_36, N85_37, I3_un3_CO1_29, 
        ADD_5x5_slow_I3_CO1_0_28, I3_un3_CO1_30, 
        ADD_5x5_slow_I3_CO1_0_29, I1_un2_CO1_13, N85_38, I3_un3_CO1_31, 
        ADD_5x5_slow_I3_CO1_0_30, I2_un4_CO1_9, 
        ADD_4x4_slow_I2_un1_CO1_0_7, N83_16, \mult1_un96_sum_1[1] , 
        N85_39, \mult1_un103_sum_1[1] , N85_40, I3_un3_CO1_32, 
        ADD_5x5_slow_I3_CO1_0_31, \mult1_un89_sum_1[1] , N85_41, N89_9, 
        N83_17, N83_18, I3_un3_CO1_33, ADD_5x5_slow_I3_CO1_0_32, 
        N85_42, I2_un1_CO1_44, I2_un1_CO1_45, I2_un4_CO1_10, 
        ADD_4x4_slow_I2_un1_CO1_0_8, I2_un1_CO1_46, I2_un4_CO1_11, 
        ADD_4x4_slow_I2_un1_CO1_0_9, I2_un4_CO1_12, 
        ADD_4x4_slow_I2_un1_CO1_0_10, I2_un4_CO1_13, 
        ADD_4x4_slow_I2_un1_CO1_0_11, I2_un1_CO1_47, I2_un1_CO1_48, 
        I2_un1_CO1_1_3, I2_un4_CO1_14, I2_un4_CO1_15, 
        ADD_5x5_slow_I2_un1_CO1_0_0, I2_un1_CO1_1_4, I2_un4_CO1_16, 
        I2_un4_CO1_17, I2_un4_CO1_18, ADD_5x5_slow_I2_un1_CO1_0_1, 
        N85_1_0, I2_un4_CO1_19, I2_un1_CO1_1_5, I2_un4_CO1_20, 
        ADD_5x5_slow_I2_un1_CO1_0_2, I1_un3_CO1_4, I2_un1_CO1_1_6, 
        I2_un1_CO1_1_7, ADD_5x5_slow_I3_CO1_0_33, I2_un4_CO1_21, 
        I2_un4_CO1_22, ADD_5x5_slow_I2_un1_CO1_0_3, I1_un3_CO1_5, 
        ADD_4x4_slow_I2_un1_CO1_0_12, I1_un3_CO1_6, 
        ADD_5x5_slow_I3_CO1_0_tz, I2_un4_CO1_23, 
        ADD_5x5_slow_I2_un1_CO1_0_4, ADD_5x5_slow_I2_un1_CO1_0_tz, 
        N85_1_1, ADD_4x4_slow_I2_un1_CO1_0_tz, N74_1_0, I2_un1_CO1_1_8, 
        ADD_4x4_slow_I2_un1_CO1_0_tz_0, I1_un3_CO1_7, I2_un1_CO1_1_9, 
        N74_1_1, ADD_5x5_slow_I3_CO1_0_34, ADD_5x5_slow_I3_CO1_0_tz_0, 
        ADD_5x5_slow_I2_un1_CO1_0_5, I1_un3_CO1_8, I2_un1_CO1_1_10, 
        I2_un4_CO1_24, ADD_5x5_slow_I2_un1_CO1_0_6, I1_un3_CO1_9, 
        I2_un1_CO1_1_11, N74_1_2, I2_un4_CO1_25, 
        ADD_5x5_slow_I2_un1_CO1_0_7, N85_1_2, ADD_5x5_slow_I3_CO1_0_35, 
        I2_un4_CO1_26, I2_un1_CO1_1_12, N74_1_3, 
        ADD_5x5_slow_I3_CO1_0_tz_1, ADD_4x4_slow_I2_un1_CO1_0_13, 
        ADD_4x4_slow_I2_un1_CO1_0_tz_1, ADD_5x5_slow_I2_un1_CO1_0_8, 
        ADD_5x5_slow_I2_un1_CO1_0_tz_0, ADD_4x4_slow_I2_un1_CO1_0_14, 
        I2_un4_CO1_27, N74_1_4, ADD_5x5_slow_I2_un1_CO1_0_9, 
        ADD_5x5_slow_I2_un1_CO1_0_tz_1, I1_un3_CO1_10, N74_1_5, 
        I2_un1_CO1_1_13, I2_un1_CO1_1_14, I2_un4_CO1_28, N74_1_6, 
        ADD_5x5_slow_I2_un1_CO1_0_10, N74_1_7, I2_un4_CO1_29, 
        ADD_5x5_slow_I2_un1_CO1_0_11, ADD_5x5_slow_I2_un1_CO1_0_12, 
        I1_un3_CO1_11, N74_1_8, ADD_5x5_slow_I3_CO1_0_36, 
        I2_un1_CO1_1_15, I2_un4_CO1_30, N74_1_9, 
        ADD_5x5_slow_I2_un1_CO1_0_13, I1_un3_CO1_12, 
        ADD_4x4_slow_I2_un1_CO1_0_15, ADD_4x4_slow_I2_un1_CO1_0_tz_2, 
        I2_un4_CO1_31, ADD_5x5_slow_I2_un1_CO1_0_14, 
        ADD_4x4_slow_I2_un1_CO1_0_16, I1_un3_CO1_13, I2_un1_CO1_1_tz_0, 
        I2_un1_CO1_1_tz_1, I2_un1_CO1_1_tz_2, I2_un1_CO1_1_tz_3, 
        I2_un1_CO1_1_tz_4, I3_un3_CO1_34, I2_un4_CO1_32, I2_un1_CO1_49, 
        I3_un3_CO1_35, I3_un3_CO1_36, I2_un5_CO1_2, I2_un5_CO1_3, 
        \d2_RNO_0[0]_net_1 , \d2_RNO[0]_net_1 , \d4_RNO_0[1]_net_1 , 
        \d4_RNO[1]_net_1 , \d8_RNO_0[2]_net_1 , \d8_RNO[2]_net_1 , 
        I1_un5_CO1_3, \rd_RNO[0]_net_1 , I1_un3_CO1_14, I2_un5_CO1_4, 
        I2_un5_CO1_5, I2_un5_CO1_6, I2_un5_CO1_7, I1_un2_CO1_14, 
        \d6_RNO[2]_net_1 , I_14_4, \d7_RNO[2]_net_1 , I_14_3, 
        \d6_RNO[1]_net_1 , \DWACT_ADD_CI_0_partial_sum[1] , 
        \d7_RNO[1]_net_1 , I_12_3, \d6_RNO[0]_net_1 , 
        \d7_RNO[0]_net_1 , \DWACT_ADD_CI_0_partial_sum[0] , 
        \d5_RNO[2]_net_1 , I_14_5, \d5_RNO[1]_net_1 , I_12_4, 
        \d5_RNO[0]_net_1 , \DWACT_ADD_CI_0_partial_sum_0[0] , 
        \d3_RNO[1]_net_1 , I_10, \d3_RNO[0]_net_1 , 
        \DWACT_ADD_CI_0_partial_sum_1[0] , \d7_RNO_0[1]_net_1 , 
        \d7_RNO_0[0]_net_1 , \d5_RNO_0[2]_net_1 , \d7_RNO_0[2]_net_1 , 
        \d5_RNO_0[1]_net_1 , \d6_RNO_0[1]_net_1 , \d5_RNO_0[0]_net_1 , 
        \d6_RNO_0[2]_net_1 , \d3_RNO_0[1]_net_1 , \d3_RNO_0[0]_net_1 , 
        \d6_RNO_0[0]_net_1 , \d2[0]_net_1 , \d4[1]_net_1 , 
        \d8[2]_net_1 , \d3[0]_net_1 , \d5[0]_net_1 , \d6[0]_net_1 , 
        \d7[0]_net_1 , \d3[1]_net_1 , \d5[1]_net_1 , \d6[1]_net_1 , 
        \d7[1]_net_1 , \d5[2]_net_1 , \d6[2]_net_1 , \d7[2]_net_1 , 
        \DWACT_ADD_CI_0_g_array_1_0[0] , 
        \DWACT_ADD_CI_0_pog_array_0[0] , \DWACT_ADD_CI_0_TMP_0[0] , 
        \DWACT_ADD_CI_0_g_array_0_1[0] , 
        \DWACT_ADD_CI_0_partial_sum[2] , 
        \DWACT_ADD_CI_0_partial_sum_0[1] , 
        \DWACT_ADD_CI_0_partial_sum_0[2] , 
        \DWACT_ADD_CI_0_g_array_0_1_0[0] , 
        \DWACT_ADD_CI_0_partial_sum_1[2] , 
        \DWACT_ADD_CI_0_partial_sum_1[1] , \DWACT_ADD_CI_0_TMP_1[0] , 
        GND, VCC;
    
    XOR2 \un2_d6_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_12), .B(N83_10), .Y(
        \mult1_un75_sum_0[3] ));
    XNOR2 \un2_d5_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un54_sum_0[2] ), .B(\mult1_un54_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_24));
    OA1 
        \un2_d7_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(N85_11), .B(\mult1_un40_sum[4] ), .C(\mult1_un40_sum_0[1] )
        , .Y(I2_un1_CO1_1_14));
    XOR2 \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_0_2), .B(N85_21), .Y(\mult1_un159_sum[2] )
        );
    XOR2 \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I2_S_0  
        (.A(\mult1_un166_sum[1] ), .B(\mult1_un166_sum_0[4] ), .Y(
        ADD_5x5_slow_I2_S_0_1));
    XOR2 \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I4_Y  (
        .A(N89), .B(ADD_5x5_slow_I4_Y_2_0), .Y(\mult1_un89_sum[4] ));
    XOR2 \un2_d3_if_generate_plus.mult1_un1_sum_I_7  (.A(
        ADD_4x4_slow_I1_S), .B(ADD_4x4_slow_I3_Y), .Y(
        \DWACT_ADD_CI_0_partial_sum_1[1] ));
    XNOR3 
        \un2_d7_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_9), .B(ADD_5x5_slow_I4_Y_0_6), .C(
        \mult1_un138_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_8));
    AO1 
        \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N85_4), .B(\mult1_un82_sum_0[4] ), .C(I2_un1_CO1_1_11), .Y(
        I2_un1_CO1_23));
    XNOR2 \un2_d3_if_generate_plus.mult1_un40_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[19]_net_1 ), .B(\rd[20]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_17));
    NOR2 \d7_RNO[0]  (.A(reset_c), .B(\DWACT_ADD_CI_0_partial_sum[0] ), 
        .Y(\d7_RNO[0]_net_1 ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_14), .B(\mult1_un124_sum_0[2] ), .Y(
        I3_un3_CO1_8));
    NOR3B 
        \un2_d5_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I2_un5_CO1  
        (.A(\rd[5]_net_1 ), .B(\mult1_un131_sum_0[4] ), .C(
        \rd[6]_net_1 ), .Y(I2_un5_CO1_7));
    AX1D \un2_d3_if_generate_plus.mult1_un173_sum_ADD_4x4_slow_I3_Y_1  
        (.A(I1_un2_CO1_0), .B(ADD_4x4_slow_I1_CO1_0), .C(
        ADD_4x4_slow_I3_Y_0), .Y(ADD_4x4_slow_I3_Y_1));
    MAJ3 
        \un2_d7_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\mult1_un61_sum[4] ), .B(N85_6), .C(\mult1_un61_sum_0[1] ), 
        .Y(I2_un1_CO1_29));
    XNOR3 
        \un2_d5_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_20), .B(ADD_5x5_slow_I4_Y_0_15), .C(
        \mult1_un110_sum_0[4] ), .Y(ADD_5x5_slow_I4_Y_2_19));
    AX1D \un2_d3_if_generate_plus.mult1_un54_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_13), .B(ADD_4x4_slow_I2_un1_CO1_0_11), .C(
        ADD_4x4_slow_I3_Y_2_15), .Y(\mult1_un54_sum[3] ));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_15), .B(\mult1_un110_sum[2] ), .Y(I3_un3_CO1_19)
        );
    AX1D \un2_d7_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_21), .B(ADD_5x5_slow_I3_CO1_0_20), .C(
        ADD_5x5_slow_I4_Y_2_18), .Y(\mult1_un110_sum[4] ));
    XNOR3 \un2_d7_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I2_S  (
        .A(N85_10), .B(ADD_4x4_slow_I1_S_0_19), .C(\mult1_un26_sum[4] )
        , .Y(\mult1_un33_sum[2] ));
    DFN1C0 \rd[3]  (.D(\rd[2]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[3]_net_1 ));
    NOR2 \d7_RNO[2]  (.A(reset_c), .B(I_14_3), .Y(\d7_RNO[2]_net_1 ));
    XNOR2 
        \un2_d7_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_4), .B(\mult1_un103_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_18));
    XOR3 \un2_d7_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un68_sum[4] ), .B(\mult1_un68_sum_0[1] ), .C(N85_5), 
        .Y(\mult1_un75_sum[2] ));
    AO13 \un2_d5_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I3_CO1  
        (.A(I2_un1_CO1_30), .B(\mult1_un61_sum_0[2] ), .C(
        \mult1_un61_sum_0[4] ), .Y(N89_7));
    XNOR2 \un2_d7_if_generate_plus.mult1_un1_sum_I_9  (.A(
        ADD_5x5_slow_I4_Y_0_27), .B(\rd[0]_net_1 ), .Y(
        \DWACT_ADD_CI_0_partial_sum[0] ));
    NOR2B 
        \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(N74_0), .B(\mult1_un152_sum_0[1] ), .Y(I2_un4_CO1_6));
    AOI1B 
        \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I1_CO1_0  
        (.A(\mult1_un145_sum[4] ), .B(\rd[4]_net_1 ), .C(\rd[3]_net_1 )
        , .Y(ADD_5x5_slow_I1_CO1_0));
    XNOR2 
        \un2_d5_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un124_sum_0[2] ), .B(\mult1_un124_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_11));
    OR2 
        \un2_d5_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(ADD_5x5_slow_I2_un1_CO1_0_13), .B(I2_un4_CO1_30), .Y(
        I2_un1_CO1_39));
    XNOR3 
        \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_10), .B(ADD_5x5_slow_I4_Y_0_7), .C(
        \mult1_un145_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_9));
    XOR2 \un2_d6_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_10), .B(\mult1_un89_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_8));
    XNOR2 
        \un2_d6_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_8), .B(\mult1_un96_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_8));
    AO1 
        \un2_d3_if_generate_plus.mult1_un96_sum_ADD_4x4_slow_I2_un1_CO1  
        (.A(N74_9), .B(\mult1_un89_sum[1] ), .C(
        ADD_4x4_slow_I2_un1_CO1_0_14), .Y(I2_un1_CO1_44));
    XNOR2 
        \un2_d5_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un117_sum_0[2] ), .B(\mult1_un117_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_13));
    OR2 
        \un2_d5_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(ADD_5x5_slow_I2_un1_CO1_0_7), .B(I2_un4_CO1_25), .Y(
        I2_un1_CO1_25));
    OR2A 
        \un2_d5_if_generate_plus.mult1_un19_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(\rd[23]_net_1 ), .B(I1_un3_CO1), .Y(
        ADD_5x5_slow_I2_un1_CO1_0));
    XNOR3 \un2_d5_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un40_sum_0[4] ), .B(\mult1_un40_sum_0[2] ), .C(
        I2_un1_CO1_35), .Y(ADD_5x5_slow_I4_Y_1_11));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un110_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[9]_net_1 ), .B(\rd[10]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_7));
    XNOR2 \un2_d6_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_18), .B(I2_un4_CO1_0), .Y(
        ADD_5x5_slow_I2_S_1_16));
    XOR3 \un2_d7_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un89_sum[4] ), .B(\mult1_un89_sum_0[1] ), .C(N85_8), 
        .Y(\mult1_un96_sum[2] ));
    XNOR2 \un2_d7_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un61_sum[2] ), .B(\mult1_un61_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_23));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_25), .B(\mult1_un82_sum_0[2] ), .C(
        \mult1_un82_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_32));
    XOR3 \un2_d5_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un82_sum[4] ), .B(\mult1_un82_sum_1[1] ), .C(N85_42), 
        .Y(\mult1_un89_sum_0[2] ));
    XNOR2 \un2_d3_if_generate_plus.mult1_un33_sum_ADD_4x4_slow_I3_Y_2  
        (.A(ADD_4x4_slow_I3_Y_1_10), .B(\mult1_un26_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_2_18));
    AX1D \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_28), .B(ADD_5x5_slow_I3_CO1_0_27), .C(
        ADD_5x5_slow_I4_Y_2_9), .Y(\mult1_un152_sum_0[4] ));
    XNOR2 \un2_d6_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_13), .B(\mult1_un61_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_13));
    XNOR3 \un2_d3_if_generate_plus.mult1_un61_sum_ADD_4x4_slow_I3_Y_2  
        (.A(N74_15), .B(ADD_4x4_slow_I3_Y_0_9), .C(\mult1_un54_sum[3] )
        , .Y(ADD_4x4_slow_I3_Y_2_14));
    OR2 
        \un2_d7_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N85), .B(\mult1_un19_sum[1] ), .Y(I2_un1_CO1_0));
    AO13 
        \un2_d3_if_generate_plus.mult1_un131_sum_ADD_4x4_slow_I2_un1_CO1  
        (.A(N74_4), .B(\mult1_un124_sum[1] ), .C(\mult1_un124_sum[3] ), 
        .Y(I2_un1_CO1_46));
    XNOR2 
        \un2_d7_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un124_sum[2] ), .B(\mult1_un124_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_8));
    AO18 \un2_d5_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un68_sum_0[4] ), .B(\rd[14]_net_1 ), .C(
        \rd[15]_net_1 ), .Y(N85_30));
    NOR2A \un2_d3_if_generate_plus.mult1_un1_sum_I_1  (.A(
        ADD_4x4_slow_I3_Y), .B(\rd[0]_net_1 ), .Y(
        \DWACT_ADD_CI_0_TMP_1[0] ));
    OR3 \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I1_CO1  (
        .A(I1_un5_CO1), .B(I1_un3_CO1_0), .C(I1_un2_CO1_2), .Y(N85_4));
    DFN1E1 \cur_rand_1[9]  (.D(\d2[0]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[9]));
    NOR2A \d5_RNO_0[0]  (.A(\DWACT_ADD_CI_0_partial_sum_0[0] ), .B(
        reset_c), .Y(\d5_RNO_0[0]_net_1 ));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_2), .B(\mult1_un54_sum_0[2] ), .C(
        \mult1_un54_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_23));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un173_sum_ADD_4x4_slow_I3_Y_0  
        (.A(\mult1_un159_sum_0[1] ), .B(\mult1_un159_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_0));
    XNOR2 
        \un2_d7_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un117_sum[2] ), .B(\mult1_un117_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_10));
    DFN1C0 \rd[19]  (.D(\rd[18]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[19]_net_1 ));
    OA1 
        \un2_d5_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(I1_un3_CO1_5), .B(\mult1_un124_sum_0[1] ), .C(
        \mult1_un124_sum_0[4] ), .Y(ADD_5x5_slow_I2_un1_CO1_0_3));
    XOR2 \un2_d7_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_0_0), .B(N85_18), .Y(\mult1_un166_sum[2] )
        );
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_35), .B(\mult1_un40_sum_0[2] ), .Y(
        I3_un3_CO1_23));
    AO1 \un2_d3_if_generate_plus.mult1_un110_sum_ADD_4x4_slow_I1_CO1  
        (.A(\mult1_un103_sum[3] ), .B(\rd[9]_net_1 ), .C(N74_1_3), .Y(
        N74_7));
    XOR3 \un2_d7_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un40_sum[4] ), .B(\mult1_un40_sum_0[1] ), .C(N85_11), 
        .Y(\mult1_un47_sum[2] ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(\mult1_un40_sum_1[1] ), .B(N85_28), .Y(I2_un4_CO1_28));
    DFN1C0 \rd[22]  (.D(\rd[21]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[22]_net_1 ));
    AO13 \un2_d7_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I3_CO1  
        (.A(I2_un1_CO1_32), .B(\mult1_un47_sum[2] ), .C(
        \mult1_un47_sum[4] ), .Y(N89_4));
    XOR3 \un2_d7_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un33_sum[4] ), .B(\mult1_un33_sum_0[1] ), .C(N85_14), 
        .Y(\mult1_un40_sum[2] ));
    XNOR2 \un2_d5_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_16), .B(\mult1_un19_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_41));
    OR2 
        \un2_d5_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I2_un1_CO1_0_tz  
        (.A(\mult1_un61_sum_1[1] ), .B(I1_un3_CO1_10), .Y(
        ADD_5x5_slow_I2_un1_CO1_0_tz_1));
    XNOR2 \un2_d7_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I2_S  (
        .A(N85), .B(\mult1_un19_sum[1] ), .Y(\mult1_un26_sum[2] ));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un152_sum_ADD_4x4_slow_I1_un2_CO1  
        (.A(\mult1_un145_sum[3] ), .B(\rd[4]_net_1 ), .Y(I1_un2_CO1_4));
    NOR2 \d6_RNO[0]  (.A(reset_c), .B(\rd[0]_net_1 ), .Y(
        \d6_RNO[0]_net_1 ));
    XOR3 \un2_d5_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un159_sum_0[4] ), .B(\mult1_un159_sum_1[1] ), .C(
        N85_20), .Y(\mult1_un166_sum_1[2] ));
    AO1 
        \un2_d5_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N85_34), .B(\mult1_un33_sum_1[1] ), .C(
        ADD_5x5_slow_I2_un1_CO1_0_12), .Y(I2_un1_CO1_37));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un110_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(N74_1_3), .B(\mult1_un103_sum_0[1] ), .C(
        \mult1_un103_sum[3] ), .Y(ADD_4x4_slow_I2_un1_CO1_0_8));
    AO1 
        \un2_d5_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N85_39), .B(\mult1_un96_sum_1[1] ), .C(
        ADD_5x5_slow_I2_un1_CO1_0_5), .Y(I2_un1_CO1_22));
    XOR2 \un2_d7_if_generate_plus.mult1_un1_sum_I_10  (.A(
        ADD_5x5_slow_I2_S_0_11), .B(ADD_5x5_slow_I4_Y_0_27), .Y(
        \DWACT_ADD_CI_0_partial_sum[2] ));
    AO1 \un2_d3_if_generate_plus.mult1_un89_sum_ADD_4x4_slow_I1_CO1  (
        .A(\mult1_un82_sum[3] ), .B(\rd[12]_net_1 ), .C(N74_1_4), .Y(
        N74_10));
    XOR2 \un2_d3_if_generate_plus.mult1_un117_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_6), .B(\mult1_un110_sum[3] ), .Y(
        \mult1_un117_sum[1] ));
    XOR2 \un2_d6_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_3), .B(\mult1_un138_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_1));
    XOR2 \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I3_Y_1  
        (.A(ADD_4x4_slow_I3_Y_0_1), .B(N74_1), .Y(
        ADD_4x4_slow_I3_Y_1_0));
    OR2 
        \un2_d5_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(ADD_5x5_slow_I2_un1_CO1_0_6), .B(I2_un4_CO1_24), .Y(
        I2_un1_CO1_24));
    AX1D \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I4_Y_1  
        (.A(I2_un1_CO1_1_1), .B(I2_un5_CO1_0), .C(
        ADD_5x5_slow_I4_Y_0_22), .Y(ADD_5x5_slow_I4_Y_1_0));
    XNOR2 
        \un2_d7_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_2), .B(\mult1_un110_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_16));
    XNOR2 \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un68_sum[2] ), .B(\mult1_un68_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_21));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(\mult1_un26_sum[4] ), .B(N85_10), .C(
        ADD_4x4_slow_I1_S_0_19), .Y(I2_un1_CO1_1_15));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I2_un5_CO1  
        (.A(I1_un3_CO1_14), .B(\mult1_un68_sum_0[4] ), .Y(I2_un5_CO1_0)
        );
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(\mult1_un33_sum_0[1] ), .B(N85_14), .Y(I2_un4_CO1_29));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un89_sum_ADD_4x4_slow_I1_un3_CO1  
        (.A(\rd[12]_net_1 ), .B(\rd[13]_net_1 ), .Y(I1_un3_CO1_0));
    XNOR2 \un2_d7_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_9), .B(\mult1_un54_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_31));
    DFN1P1C1 \d7[2]  (.D(I_14_3), .CLK(ref_signal_c), .PRE(
        \d7_RNO_0[2]_net_1 ), .CLR(\d7_RNO[2]_net_1 ), .Q(
        \d7[2]_net_1 ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(N85_16), .B(\mult1_un124_sum_0[1] ), .Y(I2_un4_CO1_22));
    DFN1P1C1 \d3[0]  (.D(\DWACT_ADD_CI_0_partial_sum_1[0] ), .CLK(
        ref_signal_c), .PRE(\d3_RNO_0[0]_net_1 ), .CLR(
        \d3_RNO[0]_net_1 ), .Q(\d3[0]_net_1 ));
    XNOR3 
        \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I3_Y_0  
        (.A(\mult1_un138_sum[3] ), .B(ADD_4x4_slow_I1_S_0_0), .C(
        \mult1_un145_sum[3] ), .Y(ADD_4x4_slow_I3_Y_0_1));
    XA1 
        \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I1_un5_CO1  
        (.A(I2_un1_CO1_18), .B(ADD_4x4_slow_I3_Y_2_0), .C(
        \rd[2]_net_1 ), .Y(I1_un5_CO1_3));
    XNOR2 
        \un2_d5_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un152_sum_0[2] ), .B(\mult1_un152_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_3));
    XOR2 \un2_d3_if_generate_plus.mult1_un19_sum_ADD_4x4_slow_I1_S  (
        .A(\rd[22]_net_1 ), .B(\rd[23]_net_1 ), .Y(
        \mult1_un19_sum_0[1] ));
    DFN1E1 \cur_rand_1[10]  (.D(\d4[1]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[10]));
    XNOR2 \un2_d5_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_14), .B(\mult1_un54_sum_0[4] ), .Y(
        \mult1_un61_sum_1[1] ));
    DFN1P1C1 \d5[1]  (.D(I_12_4), .CLK(ref_signal_c), .PRE(
        \d5_RNO_0[1]_net_1 ), .CLR(\d5_RNO[1]_net_1 ), .Q(
        \d5[1]_net_1 ));
    AO1 
        \un2_d7_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N85_15), .B(\mult1_un131_sum[4] ), .C(I2_un1_CO1_1_5), .Y(
        I2_un1_CO1_9));
    AX1D \un2_d5_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_20), .B(ADD_5x5_slow_I3_CO1_0_19), .C(
        ADD_5x5_slow_I4_Y_2_21), .Y(\mult1_un110_sum_0[4] ));
    AND2 \un2_d7_if_generate_plus.mult1_un1_sum_I_5  (.A(
        ADD_5x5_slow_I1_S_1), .B(ADD_5x5_slow_I4_Y_0_27), .Y(
        \DWACT_ADD_CI_0_g_array_0_1[0] ));
    AO1 
        \un2_d7_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N85_10), .B(\mult1_un26_sum[4] ), .C(I2_un1_CO1_1_15), .Y(
        I2_un1_CO1_38));
    XNOR2 
        \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un159_sum_0[2] ), .B(\mult1_un159_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_1));
    XNOR2 \un2_d3_if_generate_plus.mult1_un61_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[16]_net_1 ), .B(\rd[17]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_14));
    NOR2A 
        \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I1_un3_CO1  
        (.A(\rd[13]_net_1 ), .B(\rd[14]_net_1 ), .Y(I1_un3_CO1_1));
    XOR2 \un2_d6_if_generate_plus.mult1_un1_sum_I_14  (.A(
        \DWACT_ADD_CI_0_partial_sum_0[2] ), .B(
        \DWACT_ADD_CI_0_g_array_0_1_0[0] ), .Y(I_14_4));
    AO1 
        \un2_d7_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N85_25), .B(\mult1_un103_sum[4] ), .C(I2_un1_CO1_1_8), .Y(
        I2_un1_CO1_17));
    XOR2 \un2_d6_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_15), .B(N83_11), .Y(
        \mult1_un54_sum_0[3] ));
    AOI1B 
        \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_CO1_0  
        (.A(\mult1_un166_sum_0[4] ), .B(\rd[1]_net_1 ), .C(
        \rd[0]_net_1 ), .Y(ADD_5x5_slow_I1_CO1_0_2));
    OR2 
        \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(I2_un5_CO1_5), .B(I2_un1_CO1_1_12), .Y(I2_un1_CO1_27));
    AO13 \un2_d7_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un89_sum[4] ), .B(\rd[11]_net_1 ), .C(
        \rd[12]_net_1 ), .Y(N85_8));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_22), .B(\mult1_un96_sum_0[2] ), .Y(
        I3_un3_CO1_34));
    AX1D \un2_d7_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_12), .B(ADD_5x5_slow_I3_CO1_0_11), .C(
        ADD_5x5_slow_I4_Y_2_2), .Y(\mult1_un166_sum[4] ));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_5), .B(\mult1_un131_sum[2] ), .C(
        \mult1_un131_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_16));
    MAJ3 
        \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\mult1_un75_sum_0[4] ), .B(N85_3), .C(\mult1_un75_sum[1] ), 
        .Y(I2_un1_CO1_26));
    OR2 \un2_d7_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I3_CO1  
        (.A(ADD_5x5_slow_I3_CO1_0_33), .B(I3_un3_CO1_35), .Y(N89_5));
    AO13 
        \un2_d3_if_generate_plus.mult1_un68_sum_ADD_4x4_slow_I2_un1_CO1  
        (.A(N74_13), .B(\mult1_un61_sum[1] ), .C(\mult1_un61_sum[3] ), 
        .Y(I2_un1_CO1_43));
    XOR2 \un2_d7_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_0_3), .B(N85_23), .Y(\mult1_un145_sum[2] )
        );
    DFN1P1C1 \d7[1]  (.D(I_12_3), .CLK(ref_signal_c), .PRE(
        \d7_RNO_0[1]_net_1 ), .CLR(\d7_RNO[1]_net_1 ), .Q(
        \d7[1]_net_1 ));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_7), .B(\mult1_un138_sum[2] ), .Y(I3_un3_CO1_18));
    AX1D \un2_d7_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_3), .B(ADD_5x5_slow_I3_CO1_0_2), .C(
        ADD_5x5_slow_I4_Y_2_29), .Y(\mult1_un68_sum[4] ));
    AX1D \un2_d5_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_30), .B(ADD_5x5_slow_I3_CO1_0_29), .C(
        ADD_5x5_slow_I4_Y_2_5), .Y(\mult1_un166_sum_0[4] ));
    AO1A \un2_d5_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un152_sum_0[4] ), .B(\rd[2]_net_1 ), .C(N85_1_0), 
        .Y(N85_36));
    XNOR3 
        \un2_d3_if_generate_plus.mult1_un166_sum_ADD_4x4_slow_I3_Y_2  
        (.A(N74_0), .B(ADD_4x4_slow_I3_Y_0_0), .C(\mult1_un159_sum[3] )
        , .Y(ADD_4x4_slow_I3_Y_2));
    AO18 \un2_d5_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un40_sum_0[4] ), .B(\rd[18]_net_1 ), .C(
        \rd[19]_net_1 ), .Y(N85_28));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(\mult1_un75_sum_0[1] ), .B(I2_un1_CO1_1_tz_3), .Y(
        I2_un1_CO1_1_12));
    AO13 \un2_d6_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un124_sum_0[3] ), .B(\rd[7]_net_1 ), .C(
        \rd[8]_net_1 ), .Y(N83_5));
    XOR2 \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_11), .B(\mult1_un75_sum_0[4] ), .Y(
        \mult1_un82_sum[1] ));
    XOR2 \un2_d3_if_generate_plus.mult1_un33_sum_ADD_4x4_slow_I3_Y  (
        .A(ADD_4x4_slow_I3_Y_2_18), .B(I2_un1_CO1_48), .Y(
        \mult1_un33_sum[3] ));
    AO1 
        \un2_d7_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I3_CO1_0_tz  
        (.A(\mult1_un110_sum[1] ), .B(N85_26), .C(\mult1_un110_sum[2] )
        , .Y(ADD_5x5_slow_I3_CO1_0_tz));
    MAJ3 
        \un2_d5_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\mult1_un159_sum_0[4] ), .B(N85_20), .C(
        \mult1_un159_sum_1[1] ), .Y(I2_un1_CO1_4));
    AO13 \un2_d6_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un40_sum_1[4] ), .B(\rd[19]_net_1 ), .C(
        \rd[20]_net_1 ), .Y(N83_1));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(\mult1_un117_sum_0[4] ), .B(ADD_5x5_slow_I2_un1_CO1_0_tz), 
        .Y(ADD_5x5_slow_I2_un1_CO1_0_4));
    OR2 
        \un2_d5_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(ADD_5x5_slow_I2_un1_CO1_0_10), .B(I2_un4_CO1_28), .Y(
        I2_un1_CO1_35));
    XOR2 \un2_d7_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I4_Y  (
        .A(ADD_5x5_slow_I4_Y_2_14), .B(N89_5), .Y(\mult1_un124_sum[4] )
        );
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(\mult1_un138_sum[1] ), .B(N85_23), .Y(I2_un4_CO1_19));
    OA1A 
        \un2_d3_if_generate_plus.mult1_un166_sum_ADD_4x4_slow_I1_CO1_0  
        (.A(\rd[2]_net_1 ), .B(\mult1_un159_sum[3] ), .C(\rd[1]_net_1 )
        , .Y(ADD_4x4_slow_I1_CO1_0));
    XOR2 \un2_d6_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_1), .B(N83_4), .Y(\mult1_un152_sum[3] ));
    XNOR2 \un2_d3_if_generate_plus.mult1_un89_sum_ADD_4x4_slow_I3_Y_0  
        (.A(\mult1_un75_sum_1[1] ), .B(\mult1_un75_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_0_6));
    XOR2 \un2_d7_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I4_Y  (
        .A(ADD_5x5_slow_I4_Y_2_39), .B(N89_3), .Y(\mult1_un33_sum[4] ));
    XOR2 \un2_d5_if_generate_plus.mult1_un19_sum_ADD_5x5_slow_I2_S  (
        .A(\rd[23]_net_1 ), .B(N85_1), .Y(\mult1_un19_sum_0[2] ));
    XNOR3 
        \un2_d6_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I2_S_2  
        (.A(N83), .B(ADD_5x5_slow_I2_S_2_0), .C(ADD_5x5_slow_I2_S_1), 
        .Y(ADD_5x5_slow_I2_S_2));
    XNOR2 \un2_d5_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_6), .B(\mult1_un68_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_28));
    XNOR3 
        \un2_d3_if_generate_plus.mult1_un124_sum_ADD_4x4_slow_I3_Y_1  
        (.A(\mult1_un110_sum[3] ), .B(\mult1_un110_sum_0[1] ), .C(
        N74_6), .Y(ADD_4x4_slow_I3_Y_1_3));
    AX1D \un2_d5_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_22), .B(ADD_5x5_slow_I3_CO1_0_21), .C(
        ADD_5x5_slow_I4_Y_2_34), .Y(\mult1_un54_sum_0[4] ));
    OA1 
        \un2_d7_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(N85_25), .B(\mult1_un103_sum[4] ), .C(\mult1_un103_sum[1] )
        , .Y(I2_un1_CO1_1_8));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un110_sum_ADD_4x4_slow_I1_CO1_1  
        (.A(\mult1_un103_sum[3] ), .B(\rd[9]_net_1 ), .C(
        \rd[10]_net_1 ), .Y(N74_1_3));
    AO13 \un2_d7_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un40_sum[4] ), .B(\rd[18]_net_1 ), .C(
        \rd[19]_net_1 ), .Y(N85_11));
    XNOR3 \un2_d5_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un33_sum_0[4] ), .B(\mult1_un33_sum_0[2] ), .C(
        I2_un1_CO1_37), .Y(ADD_5x5_slow_I4_Y_1_13));
    AO13 \un2_d7_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un138_sum[4] ), .B(\rd[4]_net_1 ), .C(\rd[5]_net_1 )
        , .Y(N85_23));
    XOR2 \un2_d5_if_generate_plus.mult1_un1_sum_I_12  (.A(
        ADD_5x5_slow_I1_S), .B(\DWACT_ADD_CI_0_TMP[0] ), .Y(I_12_4));
    XNOR3 \un2_d3_if_generate_plus.mult1_un47_sum_ADD_4x4_slow_I3_Y_1  
        (.A(\mult1_un33_sum[3] ), .B(\mult1_un33_sum[1] ), .C(N74_17), 
        .Y(ADD_4x4_slow_I3_Y_1_8));
    NOR2A \d7_RNO_0[2]  (.A(I_14_3), .B(reset_c), .Y(
        \d7_RNO_0[2]_net_1 ));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_36), .B(\mult1_un33_sum[2] ), .Y(I3_un3_CO1_5));
    OR3 \un2_d6_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_CO1  
        (.A(I1_un5_CO1_1), .B(I1_un3_CO1_2), .C(I1_un2_CO1_11), .Y(
        N83_14));
    OR3A 
        \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I2_un1_CO1_1_tz  
        (.A(\rd[14]_net_1 ), .B(ADD_5x5_slow_I1_CO1_0_5), .C(
        \mult1_un75_sum[4] ), .Y(I2_un1_CO1_1_tz_3));
    AO1 \un2_d3_if_generate_plus.mult1_un47_sum_ADD_4x4_slow_I1_CO1  (
        .A(\mult1_un40_sum[3] ), .B(\rd[18]_net_1 ), .C(N74_1_8), .Y(
        N74_16));
    AX1D \un2_d7_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_7), .B(ADD_5x5_slow_I3_CO1_0_6), .C(
        ADD_5x5_slow_I4_Y_2_12), .Y(\mult1_un131_sum[4] ));
    MAJ3 
        \un2_d7_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\mult1_un117_sum[4] ), .B(N85_24), .C(
        \mult1_un117_sum_1[1] ), .Y(I2_un1_CO1_13));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un152_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[3]_net_1 ), .B(\rd[4]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_2));
    XNOR3 \un2_d7_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_23), .B(ADD_5x5_slow_I4_Y_0_17), .C(
        \mult1_un89_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_22));
    OR2 \un2_d7_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I3_CO1  (
        .A(ADD_5x5_slow_I3_CO1_0_36), .B(I3_un3_CO1_36), .Y(N89_3));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un166_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(I1_un3_CO1_2), .B(\mult1_un159_sum_0[1] ), .C(
        \mult1_un159_sum[3] ), .Y(ADD_4x4_slow_I2_un1_CO1_0_5));
    NOR2A 
        \un2_d5_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I1_un3_CO1  
        (.A(\rd[15]_net_1 ), .B(\rd[16]_net_1 ), .Y(I1_un3_CO1_10));
    NOR2 
        \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_un2_CO1  
        (.A(\mult1_un166_sum_0[4] ), .B(\rd[1]_net_1 ), .Y(
        I1_un2_CO1_13));
    XOR2 \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_0_1), .B(N85_35), .Y(ADD_5x5_slow_I2_S));
    DFN1E1 \cur_rand_1[21]  (.D(\d2[0]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[21]));
    OA1A 
        \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I1_CO1_0  
        (.A(\rd[14]_net_1 ), .B(\mult1_un75_sum_0[4] ), .C(
        \rd[13]_net_1 ), .Y(ADD_5x5_slow_I1_CO1_0_4));
    XOR2 \un2_d7_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I4_Y_1  
        (.A(I2_un1_CO1_0), .B(\mult1_un19_sum[2] ), .Y(
        ADD_5x5_slow_I4_Y_1));
    OA1 
        \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(N85_21), .B(\mult1_un152_sum[4] ), .C(\mult1_un152_sum[1] )
        , .Y(I2_un1_CO1_1_4));
    NOR2A 
        \un2_d6_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_un3_CO1  
        (.A(\rd[1]_net_1 ), .B(\rd[2]_net_1 ), .Y(I1_un3_CO1_2));
    XNOR2 \un2_d3_if_generate_plus.mult1_un26_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[21]_net_1 ), .B(\rd[22]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_19));
    DFN1P1C1 \d4[1]  (.D(\rd[1]_net_1 ), .CLK(ref_signal_c), .PRE(
        \d4_RNO_0[1]_net_1 ), .CLR(\d4_RNO[1]_net_1 ), .Q(
        \d4[1]_net_1 ));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un89_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(N74_1_4), .B(\mult1_un82_sum_0[1] ), .C(
        \mult1_un82_sum[3] ), .Y(ADD_4x4_slow_I2_un1_CO1_0));
    OA1 
        \un2_d5_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(I1_un3_CO1_8), .B(\mult1_un96_sum_1[1] ), .C(
        \mult1_un96_sum_0[4] ), .Y(ADD_5x5_slow_I2_un1_CO1_0_5));
    DFN1E1 \cur_rand_1[18]  (.D(\d7[0]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[18]));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(N85_33), .B(\mult1_un26_sum_0[1] ), .Y(I2_un4_CO1_30));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_21), .B(\mult1_un89_sum[2] ), .Y(I3_un3_CO1_2));
    XOR2 \un2_d3_if_generate_plus.mult1_un103_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_8), .B(\mult1_un96_sum[3] ), .Y(
        \mult1_un103_sum_0[1] ));
    DFN1C0 \rd[14]  (.D(\rd[13]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[14]_net_1 ));
    AO18 \un2_d5_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un54_sum_0[4] ), .B(\rd[16]_net_1 ), .C(
        \rd[17]_net_1 ), .Y(N85_29));
    XOR2 \un2_d7_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_5), .B(\mult1_un117_sum[4] ), .Y(
        \mult1_un124_sum_1[1] ));
    AO18 \un2_d5_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un131_sum_0[4] ), .B(\rd[5]_net_1 ), .C(
        \rd[6]_net_1 ), .Y(N85_38));
    DFN1P1C1 \d6[1]  (.D(\DWACT_ADD_CI_0_partial_sum[1] ), .CLK(
        ref_signal_c), .PRE(\d6_RNO_0[1]_net_1 ), .CLR(
        \d6_RNO[1]_net_1 ), .Q(\d6[1]_net_1 ));
    NOR2A 
        \un2_d7_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(ADD_5x5_slow_I3_CO1_0_tz), .B(\mult1_un110_sum[4] ), .Y(
        ADD_5x5_slow_I3_CO1_0_18));
    AO13 \un2_d6_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un138_sum_0[3] ), .B(\rd[5]_net_1 ), .C(
        \rd[6]_net_1 ), .Y(N83_3));
    OA1A 
        \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I2_un5_CO1  
        (.A(\rd[1]_net_1 ), .B(ADD_5x5_slow_I1_CO1_0_0), .C(
        \mult1_un166_sum[4] ), .Y(I2_un5_CO1_3));
    XOR2 \un2_d3_if_generate_plus.mult1_un138_sum_ADD_4x4_slow_I3_Y_1  
        (.A(ADD_4x4_slow_I3_Y_0_4), .B(N74_4), .Y(
        ADD_4x4_slow_I3_Y_1_1));
    XNOR3 \un2_d7_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_38), .B(ADD_5x5_slow_I4_Y_0_26), .C(
        \mult1_un33_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_37));
    XOR2 \un2_d3_if_generate_plus.mult1_un75_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_12), .B(\mult1_un68_sum[3] ), .Y(
        \mult1_un75_sum_1[1] ));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un33_sum_ADD_4x4_slow_I1_un3_CO1  
        (.A(\rd[20]_net_1 ), .B(\rd[21]_net_1 ), .Y(I1_un3_CO1_12));
    XNOR3 
        \un2_d5_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un96_sum_0[4] ), .B(\mult1_un96_sum_0[2] ), .C(
        I2_un1_CO1_22), .Y(ADD_5x5_slow_I4_Y_1_5));
    XNOR2 
        \un2_d7_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un131_sum[2] ), .B(\mult1_un131_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_6));
    XOR2 \un2_d6_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_6), .B(\mult1_un117_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_4));
    AO1A 
        \un2_d3_if_generate_plus.mult1_un89_sum_ADD_4x4_slow_I1_CO1_1  
        (.A(\rd[13]_net_1 ), .B(\mult1_un82_sum[3] ), .C(I1_un3_CO1_0), 
        .Y(N74_1_4));
    XA1 
        \un2_d6_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I1_un5_CO1  
        (.A(N83_0), .B(ADD_5x5_slow_I2_S_2_10), .C(\rd[13]_net_1 ), .Y(
        I1_un5_CO1_0));
    AX1D \un2_d5_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_8), .B(ADD_5x5_slow_I3_CO1_0_7), .C(
        ADD_5x5_slow_I4_Y_2_15), .Y(\mult1_un131_sum_0[4] ));
    XOR2 \un2_d3_if_generate_plus.mult1_un96_sum_ADD_4x4_slow_I3_Y  (
        .A(ADD_4x4_slow_I3_Y_2_9), .B(I2_un1_CO1_44), .Y(
        \mult1_un96_sum[3] ));
    OA1 
        \un2_d5_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(N85_29), .B(\mult1_un54_sum_0[4] ), .C(
        \mult1_un54_sum_1[1] ), .Y(I2_un1_CO1_1_2));
    XNOR2 \un2_d5_if_generate_plus.mult1_un1_sum_I_9  (.A(
        ADD_5x5_slow_I4_Y), .B(\rd[0]_net_1 ), .Y(
        \DWACT_ADD_CI_0_partial_sum_0[0] ));
    NOR2B 
        \un2_d3_if_generate_plus.mult1_un75_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(N74_12), .B(\mult1_un68_sum[1] ), .Y(I2_un4_CO1_2));
    OR2 
        \un2_d5_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I2_un1_CO1_1_tz  
        (.A(\mult1_un131_sum_0[4] ), .B(N85_38), .Y(I2_un1_CO1_1_tz_4));
    XOR2 \un2_d6_if_generate_plus.mult1_un1_sum_I_10  (.A(
        ADD_5x5_slow_I1_S_0), .B(I2_un1_CO1_49), .Y(
        \DWACT_ADD_CI_0_partial_sum_0[2] ));
    DFN1P1C1 \d6[0]  (.D(\rd[0]_net_1 ), .CLK(ref_signal_c), .PRE(
        \d6_RNO_0[0]_net_1 ), .CLR(\d6_RNO[0]_net_1 ), .Q(
        \d6[0]_net_1 ));
    NOR2A 
        \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I1_un2_CO1  
        (.A(\mult1_un82_sum_0[4] ), .B(\rd[13]_net_1 ), .Y(
        I1_un2_CO1_2));
    AX1D \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_31), .B(ADD_5x5_slow_I3_CO1_0_30), .C(
        ADD_5x5_slow_I4_Y_2_11), .Y(\mult1_un145_sum[4] ));
    XOR2 \un2_d7_if_generate_plus.mult1_un19_sum_ADD_5x5_slow_I1_S_0  
        (.A(\rd[23]_net_1 ), .B(\rd[22]_net_1 ), .Y(
        \mult1_un19_sum[1] ));
    OR2 \un2_d3_if_generate_plus.mult1_un152_sum_ADD_4x4_slow_I1_CO1  
        (.A(ADD_4x4_slow_I1_CO1_0_0), .B(I1_un2_CO1_4), .Y(N74_1));
    XNOR2 \un2_d3_if_generate_plus.mult1_un68_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[15]_net_1 ), .B(\rd[16]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_13));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un145_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[4]_net_1 ), .B(\rd[5]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_0));
    XOR2 \un2_d5_if_generate_plus.mult1_un1_sum_I_10  (.A(
        ADD_5x5_slow_I2_S), .B(ADD_5x5_slow_I4_Y), .Y(
        \DWACT_ADD_CI_0_partial_sum_1[2] ));
    XNOR2 \un2_d7_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_10), .B(\mult1_un47_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_33));
    XOR2 \un2_d6_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_8), .B(\mult1_un103_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_6));
    XOR2 \un2_d6_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_14), .B(N83_8), .Y(
        \mult1_un61_sum_0[3] ));
    AO1A \un2_d5_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un82_sum[4] ), .B(\rd[12]_net_1 ), .C(N85_1_2), .Y(
        N85_42));
    XNOR3 
        \un2_d5_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_16), .B(ADD_5x5_slow_I4_Y_0_13), .C(
        \mult1_un124_sum_0[4] ), .Y(ADD_5x5_slow_I4_Y_2_15));
    XNOR2 
        \un2_d6_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_6), .B(\mult1_un110_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_6));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_13), .B(\mult1_un117_sum[2] ), .Y(I3_un3_CO1_35)
        );
    XOR2 \un2_d3_if_generate_plus.mult1_un26_sum_ADD_4x4_slow_I3_Y  (
        .A(ADD_4x4_slow_I3_Y_2_19), .B(I2_un1_CO1_47), .Y(
        \mult1_un26_sum[3] ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_33), .B(\mult1_un47_sum_0[2] ), .Y(
        I3_un3_CO1_22));
    XNOR3 \un2_d7_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un33_sum[4] ), .B(\mult1_un33_sum[2] ), .C(
        I2_un1_CO1_36), .Y(ADD_5x5_slow_I4_Y_1_12));
    XOR2 \un2_d6_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_9), .B(N83_18), .Y(
        \mult1_un96_sum_0[3] ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(\mult1_un19_sum_1[1] ), .B(N85_12), .Y(I2_un4_CO1_31));
    AO18 \un2_d5_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un159_sum_0[4] ), .B(\rd[1]_net_1 ), .C(
        \rd[2]_net_1 ), .Y(N85_20));
    OR2 
        \un2_d5_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(I2_un5_CO1_7), .B(I2_un1_CO1_1_7), .Y(I2_un1_CO1_12));
    XNOR3 \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un75_sum_0[4] ), .B(\mult1_un75_sum[2] ), .C(
        I2_un1_CO1_26), .Y(ADD_5x5_slow_I4_Y_1_1));
    XNOR3 
        \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_5), .B(ADD_5x5_slow_I4_Y_0_2), .C(
        \mult1_un152_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_4));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un96_sum_ADD_4x4_slow_I1_un3_CO1  
        (.A(\rd[11]_net_1 ), .B(\rd[12]_net_1 ), .Y(I1_un3_CO1_9));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I2_un5_CO1  
        (.A(I1_un3_CO1_7), .B(\mult1_un145_sum[4] ), .Y(I2_un5_CO1_6));
    XNOR2 \un2_d3_if_generate_plus.mult1_un40_sum_ADD_4x4_slow_I3_Y_2  
        (.A(ADD_4x4_slow_I3_Y_1_9), .B(\mult1_un33_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_2_17));
    AO13 \un2_d6_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un117_sum_0[3] ), .B(\rd[8]_net_1 ), .C(
        \rd[9]_net_1 ), .Y(N83_6));
    AOI1B 
        \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I1_CO1_0  
        (.A(\mult1_un75_sum[4] ), .B(\rd[14]_net_1 ), .C(
        \rd[13]_net_1 ), .Y(ADD_5x5_slow_I1_CO1_0_5));
    AO13 \un2_d7_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un68_sum[4] ), .B(\rd[14]_net_1 ), .C(
        \rd[15]_net_1 ), .Y(N85_5));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_14), .B(\mult1_un40_sum[2] ), .C(
        \mult1_un40_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_5));
    AX1D \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I2_S  (
        .A(I1_un2_CO1_7), .B(ADD_5x5_slow_I1_CO1_0_0), .C(
        ADD_5x5_slow_I2_S_0), .Y(ADD_5x5_slow_I2_S_0_11));
    XNOR3 
        \un2_d7_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_13), .B(ADD_5x5_slow_I4_Y_0_10), .C(
        \mult1_un124_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_12));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_8), .B(\mult1_un103_sum[2] ), .C(
        \mult1_un103_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_20));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un103_sum_ADD_4x4_slow_I1_un3_CO1  
        (.A(\rd[10]_net_1 ), .B(\rd[11]_net_1 ), .Y(I1_un3_CO1_8));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_6), .B(\mult1_un152_sum_0[2] ), .Y(
        I3_un3_CO1_14));
    OA1 
        \un2_d5_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(N85_1_2), .B(\mult1_un82_sum_1[1] ), .C(
        \mult1_un82_sum[4] ), .Y(ADD_5x5_slow_I2_un1_CO1_0_7));
    AO1 \un2_d3_if_generate_plus.mult1_un54_sum_ADD_4x4_slow_I1_CO1  (
        .A(\mult1_un47_sum[3] ), .B(\rd[17]_net_1 ), .C(N74_1_7), .Y(
        N74_15));
    OA1A 
        \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I1_CO1_0  
        (.A(\rd[3]_net_1 ), .B(\mult1_un152_sum[4] ), .C(\rd[2]_net_1 )
        , .Y(ADD_5x5_slow_I1_CO1_0_3));
    XNOR3 \un2_d7_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_29), .B(ADD_5x5_slow_I4_Y_0_23), .C(
        \mult1_un68_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_27));
    OA1 
        \un2_d5_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(N85_1_0), .B(\mult1_un152_sum_1[1] ), .C(
        \mult1_un152_sum_0[4] ), .Y(ADD_5x5_slow_I2_un1_CO1_0_1));
    DFN1C0 \rd[20]  (.D(\rd[19]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[20]_net_1 ));
    AO13 \un2_d7_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un124_sum[4] ), .B(\rd[6]_net_1 ), .C(\rd[7]_net_1 )
        , .Y(N85_22));
    AO1 
        \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N85_21), .B(\mult1_un152_sum[4] ), .C(I2_un1_CO1_1_4), .Y(
        I2_un1_CO1_3));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(N85_17), .B(\mult1_un117_sum_0[1] ), .Y(I2_un4_CO1_23));
    GND GND_i (.Y(GND));
    XOR2 \un2_d5_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I4_Y  (
        .A(ADD_5x5_slow_I4_Y_2_38), .B(N89_8), .Y(
        \mult1_un40_sum_0[4] ));
    XOR3 \un2_d7_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un96_sum[4] ), .B(\mult1_un96_sum_0[1] ), .C(N85_9), 
        .Y(\mult1_un103_sum[2] ));
    OA1 
        \un2_d7_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(N85_22), .B(\mult1_un124_sum[4] ), .C(
        \mult1_un124_sum_1[1] ), .Y(I2_un1_CO1_1_6));
    XNOR3 
        \un2_d7_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un96_sum[4] ), .B(\mult1_un96_sum[2] ), .C(
        I2_un1_CO1_19), .Y(ADD_5x5_slow_I4_Y_1_4));
    NOR2A 
        \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I1_un3_CO1  
        (.A(\rd[4]_net_1 ), .B(\rd[5]_net_1 ), .Y(I1_un3_CO1_4));
    NOR2A \un2_d6_if_generate_plus.mult1_un1_sum_I_5  (.A(
        I2_un1_CO1_49), .B(\rd[1]_net_1 ), .Y(
        \DWACT_ADD_CI_0_g_array_0_1_0[0] ));
    OA1 
        \un2_d5_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_1_0), .B(I2_un5_CO1), .C(\mult1_un110_sum_0[2] )
        , .Y(I3_un3_CO1_9));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_40), .B(\mult1_un19_sum_0[2] ), .Y(
        I3_un3_CO1_27));
    XNOR2 \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I1_S  
        (.A(ADD_4x4_slow_I1_S_0_2), .B(\mult1_un145_sum[4] ), .Y(
        \mult1_un152_sum_1[1] ));
    XNOR2 \un2_d6_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_15), .B(\mult1_un47_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_15));
    XNOR3 \un2_d7_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un47_sum[4] ), .B(\mult1_un47_sum[2] ), .C(
        I2_un1_CO1_32), .Y(ADD_5x5_slow_I4_Y_1_9));
    XOR2 \un2_d5_if_generate_plus.mult1_un1_sum_I_14  (.A(
        \DWACT_ADD_CI_0_partial_sum_1[2] ), .B(
        \DWACT_ADD_CI_0_g_array_1[0] ), .Y(I_14_5));
    DFN1C0 \rd[5]  (.D(\rd[4]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[5]_net_1 ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(\mult1_un47_sum_1[1] ), .B(I2_un1_CO1_1_tz_2), .Y(
        I2_un1_CO1_1_13));
    XNOR3 
        \un2_d3_if_generate_plus.mult1_un145_sum_ADD_4x4_slow_I3_Y_2  
        (.A(N74_3), .B(ADD_4x4_slow_I3_Y_0_3), .C(\mult1_un138_sum[3] )
        , .Y(ADD_4x4_slow_I3_Y_2_2));
    XOR3 \un2_d5_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un47_sum_0[4] ), .B(\mult1_un47_sum_1[1] ), .C(
        N85_31), .Y(\mult1_un54_sum_0[2] ));
    OA1A 
        \un2_d3_if_generate_plus.mult1_un82_sum_ADD_4x4_slow_I1_CO1_0  
        (.A(\rd[14]_net_1 ), .B(\mult1_un75_sum[3] ), .C(
        \rd[13]_net_1 ), .Y(ADD_4x4_slow_I1_CO1_0_2));
    XNOR3 \un2_d3_if_generate_plus.mult1_un82_sum_ADD_4x4_slow_I3_Y_2  
        (.A(N74_12), .B(ADD_4x4_slow_I3_Y_0_7), .C(\mult1_un75_sum[3] )
        , .Y(ADD_4x4_slow_I3_Y_2_11));
    XNOR3 
        \un2_d5_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_24), .B(ADD_5x5_slow_I4_Y_0_18), .C(
        \mult1_un96_sum_0[4] ), .Y(ADD_5x5_slow_I4_Y_2_23));
    DFN1P1C1 \d6[2]  (.D(I_14_4), .CLK(ref_signal_c), .PRE(
        \d6_RNO_0[2]_net_1 ), .CLR(\d6_RNO[2]_net_1 ), .Q(
        \d6[2]_net_1 ));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un124_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(N74_1_2), .B(\mult1_un117_sum[1] ), .C(
        \mult1_un117_sum[3] ), .Y(ADD_4x4_slow_I2_un1_CO1_0_7));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_10), .B(\mult1_un89_sum[2] ), .C(
        \mult1_un89_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_1));
    NOR2B 
        \un2_d3_if_generate_plus.mult1_un82_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(N74_11), .B(\mult1_un75_sum_1[1] ), .Y(I2_un4_CO1_8));
    XNOR3 \un2_d3_if_generate_plus.mult1_un173_sum_ADD_4x4_slow_I3_Y  
        (.A(\mult1_un166_sum[3] ), .B(ADD_4x4_slow_I3_Y_1), .C(
        I2_un1_CO1_41), .Y(ADD_4x4_slow_I3_Y));
    AO13 \un2_d6_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un75_sum_0[3] ), .B(\rd[14]_net_1 ), .C(
        \rd[15]_net_1 ), .Y(N83_0));
    NOR2A 
        \un2_d6_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I1_un3_CO1  
        (.A(\rd[6]_net_1 ), .B(\rd[7]_net_1 ), .Y(I1_un3_CO1_5));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un138_sum_ADD_4x4_slow_I3_Y_0  
        (.A(\mult1_un124_sum[1] ), .B(\mult1_un124_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_0_4));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un110_sum_ADD_4x4_slow_I3_Y_2  
        (.A(ADD_4x4_slow_I3_Y_1_5), .B(\mult1_un103_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_2_7));
    NOR2 \d5_RNO[0]  (.A(reset_c), .B(
        \DWACT_ADD_CI_0_partial_sum_0[0] ), .Y(\d5_RNO[0]_net_1 ));
    XNOR2 \un2_d5_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_16), .B(\mult1_un40_sum_0[4] ), .Y(
        \mult1_un47_sum_1[1] ));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un82_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(I1_un3_CO1_1), .B(\mult1_un75_sum_1[1] ), .C(
        \mult1_un75_sum[3] ), .Y(ADD_4x4_slow_I2_un1_CO1_0_6));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_29), .B(\mult1_un33_sum[2] ), .C(
        \mult1_un33_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_4));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_19), .B(\mult1_un138_sum[2] ), .C(
        \mult1_un138_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_17));
    OR2 \un2_d3_if_generate_plus.mult1_un145_sum_ADD_4x4_slow_I1_CO1  
        (.A(ADD_4x4_slow_I1_CO1_0_1), .B(I1_un2_CO1_5), .Y(N74_2));
    XNOR2 \un2_d3_if_generate_plus.mult1_un54_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[17]_net_1 ), .B(\rd[18]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_15));
    OR2 
        \un2_d3_if_generate_plus.mult1_un33_sum_ADD_4x4_slow_I2_un1_CO1_0_tz  
        (.A(\mult1_un26_sum[1] ), .B(I1_un3_CO1_12), .Y(
        ADD_4x4_slow_I2_un1_CO1_0_tz_2));
    AX1D \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_15), .B(ADD_5x5_slow_I3_CO1_0_14), .C(
        ADD_5x5_slow_I4_Y_2_3), .Y(ADD_5x5_slow_I4_Y));
    AX1D \un2_d5_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_14), .B(ADD_5x5_slow_I3_CO1_0_13), .C(
        ADD_5x5_slow_I4_Y_2_7), .Y(\mult1_un159_sum_0[4] ));
    XOR3 \un2_d6_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I2_S_1  
        (.A(N83_0), .B(ADD_5x5_slow_I2_S_2_10), .C(
        ADD_4x4_slow_I1_S_0_11), .Y(ADD_5x5_slow_I2_S_1_9));
    XOR2 \un2_d3_if_generate_plus.mult1_un152_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_2), .B(\mult1_un145_sum[3] ), .Y(
        \mult1_un152_sum_0[1] ));
    XOR2 \un2_d6_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_17), .B(\mult1_un40_sum_1[4] ), .Y(
        ADD_5x5_slow_I2_S_1_15));
    OR2 \un2_d5_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I3_CO1  
        (.A(ADD_5x5_slow_I3_CO1_0_34), .B(I3_un3_CO1_34), .Y(N89_9));
    XNOR2 \un2_d7_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un82_sum[2] ), .B(\mult1_un82_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_17));
    XNOR2 
        \un2_d5_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un145_sum_0[2] ), .B(\mult1_un145_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_5));
    AX1D \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I2_S  (
        .A(I1_un2_CO1), .B(ADD_5x5_slow_I1_CO1_0), .C(
        ADD_5x5_slow_I2_S_0_4), .Y(\mult1_un152_sum_0[2] ));
    XNOR3 \un2_d3_if_generate_plus.mult1_un75_sum_ADD_4x4_slow_I3_Y_1  
        (.A(\mult1_un61_sum[3] ), .B(\mult1_un61_sum[1] ), .C(N74_13), 
        .Y(ADD_4x4_slow_I3_Y_1_7));
    XOR2 \un2_d7_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I2_S_0  
        (.A(\mult1_un159_sum[1] ), .B(\mult1_un159_sum[4] ), .Y(
        ADD_5x5_slow_I2_S_0_0));
    OAI1 
        \un2_d5_if_generate_plus.mult1_un19_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(ADD_5x5_slow_I2_un1_CO1_0), .B(I2_un4_CO1), .C(
        \rd[23]_net_1 ), .Y(\mult1_un19_sum[4] ));
    AO13 \un2_d3_if_generate_plus.mult1_un33_sum_ADD_4x4_slow_I1_CO1  
        (.A(\mult1_un26_sum[3] ), .B(\rd[20]_net_1 ), .C(
        \rd[21]_net_1 ), .Y(N74_18));
    NOR2 \d7_RNO[1]  (.A(reset_c), .B(I_12_3), .Y(\d7_RNO[1]_net_1 ));
    OA1A 
        \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_CO1_0  
        (.A(\rd[1]_net_1 ), .B(\mult1_un166_sum[4] ), .C(\rd[0]_net_1 )
        , .Y(ADD_5x5_slow_I1_CO1_0_0));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un124_sum_ADD_4x4_slow_I1_CO1_1  
        (.A(\mult1_un117_sum[3] ), .B(\rd[7]_net_1 ), .C(\rd[8]_net_1 )
        , .Y(N74_1_2));
    XOR2 \un2_d7_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_4), .B(\mult1_un124_sum[4] ), .Y(
        \mult1_un131_sum_0[1] ));
    AO13 \un2_d3_if_generate_plus.mult1_un131_sum_ADD_4x4_slow_I1_CO1  
        (.A(\mult1_un124_sum[3] ), .B(\rd[6]_net_1 ), .C(\rd[7]_net_1 )
        , .Y(N74_4));
    XNOR2 \un2_d6_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_11), .B(\mult1_un75_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_10));
    XNOR3 \un2_d5_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_33), .B(ADD_5x5_slow_I4_Y_0_25), .C(
        \mult1_un54_sum_0[4] ), .Y(ADD_5x5_slow_I4_Y_2_32));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_9), .B(\mult1_un131_sum[2] ), .Y(I3_un3_CO1_17));
    NOR2B 
        \un2_d3_if_generate_plus.mult1_un40_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(N74_17), .B(\mult1_un33_sum[1] ), .Y(I2_un4_CO1_11));
    XOR2 \un2_d6_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_13), .B(\mult1_un68_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_11));
    MAJ3 
        \un2_d7_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\mult1_un110_sum[4] ), .B(N85_26), .C(\mult1_un110_sum[1] )
        , .Y(I2_un1_CO1_15));
    XOR3 \un2_d5_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un96_sum_0[4] ), .B(\mult1_un96_sum_1[1] ), .C(
        N85_39), .Y(\mult1_un103_sum_0[2] ));
    XNOR3 \un2_d3_if_generate_plus.mult1_un54_sum_ADD_4x4_slow_I3_Y_2  
        (.A(N74_16), .B(ADD_4x4_slow_I3_Y_0_10), .C(
        \mult1_un47_sum[3] ), .Y(ADD_4x4_slow_I3_Y_2_15));
    DFN1E1 \cur_rand_1[17]  (.D(\d6[2]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[17]));
    NOR2 \d6_RNO[1]  (.A(reset_c), .B(\DWACT_ADD_CI_0_partial_sum[1] ), 
        .Y(\d6_RNO[1]_net_1 ));
    XNOR2 
        \un2_d6_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_2), .B(\mult1_un138_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_2));
    XNOR2 
        \un2_d6_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_4), .B(\mult1_un124_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_4));
    NOR2A \d7_RNO_0[1]  (.A(I_12_3), .B(reset_c), .Y(
        \d7_RNO_0[1]_net_1 ));
    OR2 \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_CO1  
        (.A(ADD_5x5_slow_I1_CO1_0_2), .B(I1_un2_CO1_13), .Y(N85_35));
    AO13 \un2_d3_if_generate_plus.mult1_un103_sum_ADD_4x4_slow_I1_CO1  
        (.A(\mult1_un96_sum[3] ), .B(\rd[10]_net_1 ), .C(
        \rd[11]_net_1 ), .Y(N74_8));
    XOR2 \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I2_S_0  
        (.A(\mult1_un152_sum[1] ), .B(\mult1_un152_sum[4] ), .Y(
        ADD_5x5_slow_I2_S_0_2));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_30), .B(\mult1_un26_sum_0[2] ), .C(
        \mult1_un26_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_25));
    NOR2B 
        \un2_d3_if_generate_plus.mult1_un138_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(N74_3), .B(\mult1_un131_sum[1] ), .Y(I2_un4_CO1_4));
    NOR2A 
        \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I1_un3_CO1  
        (.A(\rd[3]_net_1 ), .B(\rd[4]_net_1 ), .Y(I1_un3_CO1_7));
    XOR2 \un2_d6_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_9), .B(\mult1_un96_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_7));
    OR2 \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I1_CO1  (
        .A(ADD_5x5_slow_I1_CO1_0_4), .B(I1_un2_CO1_1), .Y(N85_3));
    XNOR3 
        \un2_d7_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_15), .B(ADD_5x5_slow_I4_Y_0_12), .C(
        \mult1_un117_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_14));
    XOR2 \un2_d7_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I4_Y  (
        .A(ADD_5x5_slow_I4_Y_2_31), .B(N89_2), .Y(\mult1_un61_sum[4] ));
    AO13 \un2_d6_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un145_sum_0[3] ), .B(\rd[4]_net_1 ), .C(
        \rd[5]_net_1 ), .Y(N83_4));
    XOR2 \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I4_Y  (
        .A(N89_0), .B(ADD_5x5_slow_I4_Y_2), .Y(\mult1_un82_sum[4] ));
    OA1 
        \un2_d7_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(N85_14), .B(\mult1_un33_sum_0[1] ), .C(\mult1_un33_sum[4] )
        , .Y(ADD_5x5_slow_I2_un1_CO1_0_11));
    XOR2 \un2_d7_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I2_S_0  
        (.A(\mult1_un110_sum[1] ), .B(\mult1_un110_sum[4] ), .Y(
        ADD_5x5_slow_I2_S_0_6));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un82_sum_ADD_4x4_slow_I1_un2_CO1  
        (.A(\mult1_un75_sum[3] ), .B(\rd[14]_net_1 ), .Y(I1_un2_CO1_3));
    NOR2B 
        \un2_d3_if_generate_plus.mult1_un54_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(N74_15), .B(\mult1_un47_sum[1] ), .Y(I2_un4_CO1_13));
    MAJ3 
        \un2_d7_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\mult1_un68_sum[4] ), .B(N85_5), .C(\mult1_un68_sum_0[1] ), 
        .Y(I2_un1_CO1_28));
    AX1D \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I2_S  (
        .A(I1_un2_CO1_10), .B(ADD_5x5_slow_I1_CO1_0_5), .C(
        ADD_5x5_slow_I2_S_0_10), .Y(\mult1_un82_sum_0[2] ));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un47_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(N74_1_8), .B(\mult1_un40_sum[1] ), .C(\mult1_un40_sum[3] ), 
        .Y(ADD_4x4_slow_I2_un1_CO1_0_10));
    XOR2 \un2_d7_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_0_7), .B(N85_25), .Y(\mult1_un110_sum[2] )
        );
    XNOR2 \un2_d5_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_9), .B(\mult1_un89_sum_0[4] ), .Y(
        \mult1_un96_sum_1[1] ));
    NOR2 \d8_RNO[2]  (.A(reset_c), .B(\rd[2]_net_1 ), .Y(
        \d8_RNO[2]_net_1 ));
    XNOR2 
        \un2_d6_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_3), .B(\mult1_un131_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_3));
    AO1 
        \un2_d5_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N85_40), .B(\mult1_un103_sum_0[4] ), .C(I2_un1_CO1_1_9), 
        .Y(I2_un1_CO1_20));
    AO13 \un2_d6_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un54_sum_0[3] ), .B(\rd[17]_net_1 ), .C(
        \rd[18]_net_1 ), .Y(N83_8));
    XNOR2 \un2_d5_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I1_S  
        (.A(ADD_4x4_slow_I1_S_0_4), .B(\mult1_un124_sum_0[4] ), .Y(
        \mult1_un131_sum_1[1] ));
    DFN1C0 \rd[16]  (.D(\rd[15]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[16]_net_1 ));
    XNOR2 \un2_d3_if_generate_plus.mult1_un1_sum_I_8  (.A(
        ADD_4x4_slow_I3_Y), .B(\rd[0]_net_1 ), .Y(
        \DWACT_ADD_CI_0_partial_sum_1[0] ));
    DFN1E1 \cur_rand_1[22]  (.D(\d4[1]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[22]));
    XOR2 \un2_d7_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I2_S_0  
        (.A(\mult1_un138_sum[1] ), .B(\mult1_un138_sum[4] ), .Y(
        ADD_5x5_slow_I2_S_0_3));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un75_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(N74_1_5), .B(\mult1_un68_sum[1] ), .C(\mult1_un68_sum[3] ), 
        .Y(ADD_4x4_slow_I2_un1_CO1_0_0));
    XOR2 \un2_d3_if_generate_plus.mult1_un110_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_7), .B(\mult1_un103_sum[3] ), .Y(
        \mult1_un110_sum_0[1] ));
    XNOR2 \un2_d6_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_9), .B(\mult1_un89_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_9));
    AX1D \un2_d5_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_32), .B(ADD_5x5_slow_I3_CO1_0_31), .C(
        ADD_5x5_slow_I4_Y_2_24), .Y(\mult1_un96_sum_0[4] ));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un61_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(N74_1_6), .B(\mult1_un54_sum[1] ), .C(\mult1_un54_sum[3] ), 
        .Y(ADD_4x4_slow_I2_un1_CO1_0_1));
    NOR2A 
        \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_un2_CO1  
        (.A(\mult1_un166_sum[4] ), .B(\rd[1]_net_1 ), .Y(I1_un2_CO1_7));
    NOR2A \d6_RNO_0[0]  (.A(\rd[0]_net_1 ), .B(reset_c), .Y(
        \d6_RNO_0[0]_net_1 ));
    DFN1E1 \cur_rand_1[7]  (.D(\d3[1]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[7]));
    XOR2 \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I2_S_0  
        (.A(\mult1_un145_sum[1] ), .B(\mult1_un145_sum[4] ), .Y(
        ADD_5x5_slow_I2_S_0_4));
    OR2 \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I3_CO1  (
        .A(I3_un3_CO1_0), .B(ADD_5x5_slow_I3_CO1_0), .Y(N89_0));
    XOR2 \un2_d3_if_generate_plus.mult1_un61_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_14), .B(\mult1_un54_sum[3] ), .Y(
        \mult1_un61_sum[1] ));
    XNOR2 \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I1_S  
        (.A(ADD_4x4_slow_I1_S_0_0), .B(\mult1_un138_sum_0[4] ), .Y(
        \mult1_un145_sum[1] ));
    AO13 \un2_d3_if_generate_plus.mult1_un68_sum_ADD_4x4_slow_I1_CO1  
        (.A(\mult1_un61_sum[3] ), .B(\rd[15]_net_1 ), .C(
        \rd[16]_net_1 ), .Y(N74_13));
    MAJ3 
        \un2_d7_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\mult1_un54_sum_0[1] ), .B(\mult1_un54_sum[4] ), .C(N85_7), 
        .Y(I2_un1_CO1_31));
    XNOR3 
        \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_12), .B(ADD_5x5_slow_I4_Y_0_9), .C(
        \mult1_un138_sum_0[4] ), .Y(ADD_5x5_slow_I4_Y_2_11));
    XNOR3 \un2_d5_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_25), .B(ADD_5x5_slow_I4_Y_0_19), .C(
        \mult1_un89_sum_0[4] ), .Y(ADD_5x5_slow_I4_Y_2_24));
    XNOR2 \un2_d5_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_19), .B(\mult1_un19_sum[4] ), .Y(
        \mult1_un26_sum_0[1] ));
    DFN1P1C1 \d7[0]  (.D(\DWACT_ADD_CI_0_partial_sum[0] ), .CLK(
        ref_signal_c), .PRE(\d7_RNO_0[0]_net_1 ), .CLR(
        \d7_RNO[0]_net_1 ), .Q(\d7[0]_net_1 ));
    AO1 
        \un2_d3_if_generate_plus.mult1_un173_sum_ADD_4x4_slow_I2_un1_CO1  
        (.A(N74_20), .B(\mult1_un166_sum_0[1] ), .C(
        ADD_4x4_slow_I2_un1_CO1_0_12), .Y(I2_un1_CO1_41));
    XNOR2 \un2_d7_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un26_sum[2] ), .B(\mult1_un26_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_26));
    DFN1C0 \rd[11]  (.D(\rd[10]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[11]_net_1 ));
    AX1D \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_13), .B(ADD_5x5_slow_I3_CO1_0_12), .C(
        ADD_5x5_slow_I4_Y_2_1), .Y(ADD_5x5_slow_I4_Y_0_27));
    XOR2 \un2_d7_if_generate_plus.mult1_un1_sum_I_11  (.A(
        ADD_5x5_slow_I1_S_1), .B(ADD_5x5_slow_I4_Y_0_27), .Y(
        \DWACT_ADD_CI_0_partial_sum_0[1] ));
    OR2 
        \un2_d5_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I2_un1_CO1_1_tz  
        (.A(\mult1_un47_sum_0[4] ), .B(N85_31), .Y(I2_un1_CO1_1_tz_2));
    XNOR2 
        \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un138_sum_0[2] ), .B(\mult1_un138_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_7));
    XA1 
        \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(\mult1_un159_sum[4] ), .B(ADD_4x4_slow_I1_S_0), .C(
        I2_un1_CO1_1_tz_1), .Y(I2_un1_CO1_1_3));
    XNOR2 \un2_d5_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_12), .B(\mult1_un68_sum_0[4] ), .Y(
        \mult1_un75_sum_0[1] ));
    DFN1C0 \rd[2]  (.D(\rd[1]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[2]_net_1 ));
    AO13 \un2_d7_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un61_sum[4] ), .B(\rd[15]_net_1 ), .C(
        \rd[16]_net_1 ), .Y(N85_6));
    XNOR3 \un2_d6_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I2_S_2  
        (.A(N83_0), .B(ADD_5x5_slow_I2_S_2_10), .C(
        ADD_5x5_slow_I2_S_1_10), .Y(ADD_5x5_slow_I2_S_2_11));
    XNOR3 
        \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_2), .B(ADD_5x5_slow_I4_Y_0), .C(
        \mult1_un166_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_1));
    AX1D \un2_d3_if_generate_plus.mult1_un166_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_7), .B(ADD_4x4_slow_I2_un1_CO1_0_5), .C(
        ADD_4x4_slow_I3_Y_2), .Y(\mult1_un166_sum[3] ));
    XOR2 \un2_d7_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_7), .B(\mult1_un103_sum[4] ), .Y(
        \mult1_un110_sum[1] ));
    AX1D \un2_d5_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_27), .B(ADD_5x5_slow_I3_CO1_0_26), .C(
        ADD_5x5_slow_I4_Y_2_41), .Y(\mult1_un26_sum_0[4] ));
    XOR2 \un2_d3_if_generate_plus.mult1_un68_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_13), .B(\mult1_un61_sum[3] ), .Y(
        \mult1_un68_sum[1] ));
    AO18 \un2_d5_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un33_sum_0[4] ), .B(\rd[19]_net_1 ), .C(
        \rd[20]_net_1 ), .Y(N85_34));
    AO13 \un2_d3_if_generate_plus.mult1_un26_sum_ADD_4x4_slow_I1_CO1  
        (.A(\mult1_un19_sum[3] ), .B(\rd[21]_net_1 ), .C(
        \rd[22]_net_1 ), .Y(N74_19));
    DFN1E1 \cur_rand_1[16]  (.D(\d6[1]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[16]));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un54_sum_ADD_4x4_slow_I1_CO1_1  
        (.A(\rd[17]_net_1 ), .B(\mult1_un47_sum[3] ), .C(
        \rd[18]_net_1 ), .Y(N74_1_7));
    NOR2A 
        \un2_d5_if_generate_plus.mult1_un19_sum_ADD_5x5_slow_I1_un3_CO1  
        (.A(\rd[22]_net_1 ), .B(\rd[23]_net_1 ), .Y(I1_un3_CO1));
    XOR2 \un2_d7_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I4_Y  (
        .A(ADD_5x5_slow_I4_Y_2_20), .B(N89_6), .Y(\mult1_un103_sum[4] )
        );
    XNOR2 \un2_d5_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_15), .B(\mult1_un47_sum_0[4] ), .Y(
        \mult1_un54_sum_1[1] ));
    XOR3 \un2_d7_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un131_sum[4] ), .B(\mult1_un131_sum_0[1] ), .C(
        N85_15), .Y(\mult1_un138_sum[2] ));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un96_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(I1_un3_CO1_9), .B(\mult1_un89_sum[1] ), .C(
        \mult1_un89_sum[3] ), .Y(ADD_4x4_slow_I2_un1_CO1_0_14));
    XOR2 \un2_d3_if_generate_plus.mult1_un96_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_9), .B(\mult1_un89_sum[3] ), .Y(
        \mult1_un96_sum[1] ));
    OR2A \un2_d7_if_generate_plus.mult1_un19_sum_ADD_5x5_slow_I1_CO1  
        (.A(\rd[23]_net_1 ), .B(\rd[22]_net_1 ), .Y(N85_0));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un40_sum_ADD_4x4_slow_I1_un3_CO1  
        (.A(\rd[19]_net_1 ), .B(\rd[20]_net_1 ), .Y(I1_un3_CO1_11));
    DFN1C0 \rd[13]  (.D(\rd[12]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[13]_net_1 ));
    DFN1E1 \cur_rand_1[13]  (.D(\d5[1]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[13]));
    XNOR2 \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un68_sum_0[2] ), .B(\mult1_un68_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_22));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un131_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[6]_net_1 ), .B(\rd[7]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_4));
    OA1A 
        \un2_d7_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I1_CO1_0  
        (.A(\rd[2]_net_1 ), .B(\mult1_un159_sum[4] ), .C(\rd[1]_net_1 )
        , .Y(ADD_5x5_slow_I1_CO1_0_1));
    XNOR2 \un2_d5_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un82_sum_0[2] ), .B(\mult1_un82_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_19));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un103_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[10]_net_1 ), .B(\rd[11]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_8));
    OA1 
        \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(N85_35), .B(\mult1_un166_sum[1] ), .C(
        \mult1_un166_sum_0[4] ), .Y(ADD_5x5_slow_I2_un1_CO1_0_0));
    AX1D \un2_d3_if_generate_plus.mult1_un40_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_11), .B(ADD_4x4_slow_I2_un1_CO1_0_9), .C(
        ADD_4x4_slow_I3_Y_2_17), .Y(\mult1_un40_sum[3] ));
    DFN1C0 \rd[8]  (.D(\rd[7]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[8]_net_1 ));
    NOR2 \d2_RNO[0]  (.A(reset_c), .B(\rd[0]_net_1 ), .Y(
        \d2_RNO[0]_net_1 ));
    XOR3 \un2_d5_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un103_sum_0[4] ), .B(\mult1_un103_sum_1[1] ), .C(
        N85_40), .Y(\mult1_un110_sum_0[2] ));
    NOR2B 
        \un2_d3_if_generate_plus.mult1_un47_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(N74_16), .B(\mult1_un40_sum[1] ), .Y(I2_un4_CO1_12));
    OA1 
        \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un4_CO1_15), .B(ADD_5x5_slow_I2_un1_CO1_0_0), .C(
        \mult1_un166_sum_1[2] ), .Y(I3_un3_CO1_15));
    AO18 \un2_d5_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un96_sum_0[4] ), .B(\rd[10]_net_1 ), .C(
        \rd[11]_net_1 ), .Y(N85_39));
    XNOR2 \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_11), .B(\mult1_un75_sum[4] ), .Y(
        \mult1_un82_sum_1[1] ));
    XOR2 \un2_d3_if_generate_plus.mult1_un26_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_19), .B(\mult1_un19_sum[3] ), .Y(
        \mult1_un26_sum[1] ));
    DFN1P1C1 \d5[0]  (.D(\DWACT_ADD_CI_0_partial_sum_0[0] ), .CLK(
        ref_signal_c), .PRE(\d5_RNO_0[0]_net_1 ), .CLR(
        \d5_RNO[0]_net_1 ), .Q(\d5[0]_net_1 ));
    AO13 \un2_d7_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un26_sum[4] ), .B(\rd[20]_net_1 ), .C(
        \rd[21]_net_1 ), .Y(N85_10));
    XOR2 \un2_d3_if_generate_plus.mult1_un131_sum_ADD_4x4_slow_I3_Y  (
        .A(ADD_4x4_slow_I3_Y_2_4), .B(I2_un1_CO1_46), .Y(
        \mult1_un131_sum[3] ));
    OR2A \un2_d3_if_generate_plus.mult1_un19_sum_ADD_4x4_slow_I1_CO1  
        (.A(\rd[23]_net_1 ), .B(\rd[22]_net_1 ), .Y(N74));
    XOR2 \un2_d7_if_generate_plus.mult1_un1_sum_I_14  (.A(
        \DWACT_ADD_CI_0_partial_sum[2] ), .B(
        \DWACT_ADD_CI_0_g_array_1_0[0] ), .Y(I_14_3));
    XOR2 \un2_d6_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_7), .B(N83_16), .Y(
        \mult1_un110_sum_0[3] ));
    AO13 \un2_d6_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un47_sum_0[3] ), .B(\rd[18]_net_1 ), .C(
        \rd[19]_net_1 ), .Y(N83_11));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[3]_net_1 ), .B(\rd[2]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_1));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_14), .B(\mult1_un159_sum[2] ), .C(
        \mult1_un159_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_11));
    XOR3 \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I1_S  (
        .A(I2_un1_CO1_18), .B(ADD_4x4_slow_I3_Y_2_0), .C(
        ADD_4x4_slow_I1_S_0_1), .Y(\mult1_un159_sum_0[1] ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_10), .B(\mult1_un138_sum_0[2] ), .Y(
        I3_un3_CO1_31));
    DFN1P1C1 \d3[1]  (.D(I_10), .CLK(ref_signal_c), .PRE(
        \d3_RNO_0[1]_net_1 ), .CLR(\d3_RNO[1]_net_1 ), .Q(
        \d3[1]_net_1 ));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(\mult1_un75_sum[1] ), .B(N85_3), .Y(I2_un4_CO1_26));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_27), .B(\mult1_un61_sum[2] ), .C(
        \mult1_un61_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_2));
    XOR3 \un2_d5_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un131_sum_0[4] ), .B(\mult1_un131_sum_1[1] ), .C(
        N85_38), .Y(\mult1_un138_sum_0[2] ));
    XNOR2 \un2_d6_if_generate_plus.mult1_un1_sum_I_11  (.A(
        I2_un1_CO1_49), .B(\rd[1]_net_1 ), .Y(
        \DWACT_ADD_CI_0_partial_sum[1] ));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(\mult1_un89_sum_0[1] ), .B(I2_un1_CO1_1_tz_0), .Y(
        I2_un1_CO1_1_10));
    XO1 
        \un2_d3_if_generate_plus.mult1_un152_sum_ADD_4x4_slow_I2_un1_CO1_0_tz  
        (.A(\mult1_un138_sum[3] ), .B(ADD_4x4_slow_I1_S_0_0), .C(
        I1_un3_CO1_7), .Y(ADD_4x4_slow_I2_un1_CO1_0_tz_0));
    XOR2 \un2_d6_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_3), .B(N83_2), .Y(
        \mult1_un138_sum_0[3] ));
    XNOR2 
        \un2_d6_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_0), .B(\mult1_un152_sum[3] ), .Y(
        ADD_5x5_slow_I2_S_2_0));
    XOR2 \un2_d6_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_14), .B(\mult1_un61_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_12));
    MAJ3 
        \un2_d7_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\mult1_un145_sum_0[4] ), .B(N85_19), .C(
        \mult1_un145_sum_0[1] ), .Y(I2_un1_CO1_5));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I1_un3_CO1  
        (.A(\rd[2]_net_1 ), .B(\rd[3]_net_1 ), .Y(I1_un3_CO1_3));
    DFN1C0 \rd[1]  (.D(\rd[0]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[1]_net_1 ));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un152_sum_ADD_4x4_slow_I3_Y_0  
        (.A(\mult1_un138_sum_1[1] ), .B(\mult1_un138_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_0_2));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(N85_37), .B(\mult1_un138_sum_0[1] ), .Y(I2_un4_CO1_20));
    XNOR2 \un2_d3_if_generate_plus.mult1_un82_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[13]_net_1 ), .B(\rd[14]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_11));
    XOR2 \un2_d5_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I4_Y  (
        .A(ADD_5x5_slow_I4_Y_2_23), .B(N89_9), .Y(
        \mult1_un103_sum_0[4] ));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un131_sum_ADD_4x4_slow_I3_Y_2  
        (.A(ADD_4x4_slow_I3_Y_1_2), .B(\mult1_un124_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_2_4));
    XOR2 \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I2_S_0  
        (.A(\mult1_un75_sum_0[1] ), .B(\mult1_un75_sum[4] ), .Y(
        ADD_5x5_slow_I2_S_0_10));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_25), .B(\mult1_un82_sum_0[2] ), .Y(
        I3_un3_CO1_33));
    NOR2 \d3_RNO[0]  (.A(reset_c), .B(
        \DWACT_ADD_CI_0_partial_sum_1[0] ), .Y(\d3_RNO[0]_net_1 ));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un173_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(I1_un3_CO1_6), .B(\mult1_un166_sum_0[1] ), .C(
        \mult1_un166_sum[3] ), .Y(ADD_4x4_slow_I2_un1_CO1_0_12));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_12), .B(\mult1_un131_sum_0[2] ), .Y(
        I3_un3_CO1_29));
    OA1 
        \un2_d3_if_generate_plus.mult1_un166_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(I1_un2_CO1_0), .B(ADD_4x4_slow_I1_CO1_0), .C(
        \mult1_un159_sum_0[1] ), .Y(I2_un4_CO1_7));
    OA1 
        \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(N85_4), .B(\mult1_un82_sum_0[4] ), .C(\mult1_un82_sum[1] ), 
        .Y(I2_un1_CO1_1_11));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_22), .B(\mult1_un124_sum_0[2] ), .C(
        \mult1_un124_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_7));
    AX1D \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I4_Y_1  
        (.A(I2_un1_CO1_1_0), .B(I2_un5_CO1), .C(ADD_5x5_slow_I4_Y_0_14)
        , .Y(ADD_5x5_slow_I4_Y_1_3));
    AO13 \un2_d6_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un152_sum[3] ), .B(\rd[3]_net_1 ), .C(\rd[4]_net_1 )
        , .Y(N83));
    XOR2 \un2_d7_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_15), .B(\mult1_un47_sum[4] ), .Y(
        \mult1_un54_sum_0[1] ));
    XOR2 \un2_d6_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_3), .B(N83_13), .Y(\mult1_un40_sum_1[4] ));
    XNOR2 \un2_d5_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I1_S  
        (.A(ADD_4x4_slow_I1_S_0_7), .B(\mult1_un103_sum_0[4] ), .Y(
        \mult1_un110_sum_1[1] ));
    XNOR3 \un2_d3_if_generate_plus.mult1_un40_sum_ADD_4x4_slow_I3_Y_1  
        (.A(\mult1_un26_sum[3] ), .B(\mult1_un26_sum[1] ), .C(N74_18), 
        .Y(ADD_4x4_slow_I3_Y_1_9));
    DFN1E1 \cur_rand_1[20]  (.D(\d7[2]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[20]));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I2_un5_CO1  
        (.A(N85_8), .B(\mult1_un89_sum[4] ), .Y(I2_un5_CO1_2));
    AO13 \un2_d6_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un61_sum_0[3] ), .B(\rd[16]_net_1 ), .C(
        \rd[17]_net_1 ), .Y(N83_9));
    OA1 
        \un2_d5_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(N85_30), .B(\mult1_un68_sum_0[4] ), .C(
        \mult1_un68_sum_1[1] ), .Y(I2_un1_CO1_1_1));
    XOR2 \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_10), .B(\mult1_un82_sum_0[4] ), .Y(
        \mult1_un89_sum_0[1] ));
    AO18 \un2_d5_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un124_sum_0[4] ), .B(\rd[6]_net_1 ), .C(
        \rd[7]_net_1 ), .Y(N85_16));
    XOR3 \un2_d5_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un33_sum_0[4] ), .B(\mult1_un33_sum_1[1] ), .C(
        N85_34), .Y(\mult1_un40_sum_0[2] ));
    XOR2 \un2_d6_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_5), .B(N83_6), .Y(
        \mult1_un124_sum_0[3] ));
    AX1D \un2_d7_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_17), .B(ADD_5x5_slow_I3_CO1_0_16), .C(
        ADD_5x5_slow_I4_Y_2_10), .Y(\mult1_un138_sum[4] ));
    OA1 
        \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(I1_un3_CO1_4), .B(\mult1_un138_sum_0[1] ), .C(
        \mult1_un138_sum_0[4] ), .Y(ADD_5x5_slow_I2_un1_CO1_0_2));
    AX1D \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_6), .B(ADD_4x4_slow_I2_un1_CO1_0_4), .C(
        ADD_4x4_slow_I3_Y_2_1), .Y(\mult1_un159_sum[3] ));
    XNOR2 \un2_d3_if_generate_plus.mult1_un96_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[12]_net_1 ), .B(\rd[11]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_9));
    AO1A 
        \un2_d3_if_generate_plus.mult1_un152_sum_ADD_4x4_slow_I2_un1_CO1  
        (.A(\mult1_un145_sum[3] ), .B(ADD_4x4_slow_I2_un1_CO1_0_tz_0), 
        .C(I2_un4_CO1_32), .Y(I2_un1_CO1_18));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_28), .B(\mult1_un40_sum_0[2] ), .C(
        \mult1_un40_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_22));
    XA1 
        \un2_d3_if_generate_plus.mult1_un152_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(\mult1_un138_sum[3] ), .B(ADD_4x4_slow_I1_S_0_0), .C(N74_1)
        , .Y(I2_un4_CO1_32));
    NOR2A \d8_RNO_0[2]  (.A(\rd[2]_net_1 ), .B(reset_c), .Y(
        \d8_RNO_0[2]_net_1 ));
    OA1A 
        \un2_d3_if_generate_plus.mult1_un152_sum_ADD_4x4_slow_I1_CO1_0  
        (.A(\rd[4]_net_1 ), .B(\mult1_un145_sum[3] ), .C(\rd[3]_net_1 )
        , .Y(ADD_4x4_slow_I1_CO1_0_0));
    OR2 \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I1_CO1  
        (.A(I1_un5_CO1_3), .B(N74_1_0), .Y(N74_0));
    OR2 
        \un2_d7_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I2_un1_CO1_1_tz  
        (.A(\mult1_un89_sum[4] ), .B(N85_8), .Y(I2_un1_CO1_1_tz_0));
    XNOR3 \un2_d3_if_generate_plus.mult1_un89_sum_ADD_4x4_slow_I3_Y_2  
        (.A(N74_11), .B(ADD_4x4_slow_I3_Y_0_6), .C(\mult1_un82_sum[3] )
        , .Y(ADD_4x4_slow_I3_Y_2_10));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un54_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(N74_1_7), .B(\mult1_un47_sum[1] ), .C(\mult1_un47_sum[3] ), 
        .Y(ADD_4x4_slow_I2_un1_CO1_0_11));
    XNOR2 \un2_d5_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I1_S  
        (.A(ADD_4x4_slow_I1_S_0_1), .B(\mult1_un152_sum_0[4] ), .Y(
        \mult1_un159_sum_1[1] ));
    XOR3 \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un117_sum_0[4] ), .B(\mult1_un117_sum_0[1] ), .C(
        N85_17), .Y(\mult1_un124_sum_0[2] ));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_15), .B(\mult1_un166_sum_1[2] ), .C(
        \mult1_un166_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_14));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_20), .B(\mult1_un138_sum_0[2] ), .C(
        \mult1_un138_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_30));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_5), .B(\mult1_un145_sum[2] ), .Y(I3_un3_CO1_16));
    XOR2 \un2_d6_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_8), .B(N83_17), .Y(
        \mult1_un103_sum_0[3] ));
    AO13 \un2_d7_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un103_sum[4] ), .B(\rd[9]_net_1 ), .C(
        \rd[10]_net_1 ), .Y(N85_25));
    OR2B 
        \un2_d3_if_generate_plus.mult1_un19_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(\rd[23]_net_1 ), .B(N74), .Y(\mult1_un19_sum[3] ));
    NOR2 \d5_RNO[2]  (.A(reset_c), .B(I_14_5), .Y(\d5_RNO[2]_net_1 ));
    XOR2 \un2_d6_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_16), .B(N83_1), .Y(
        \mult1_un47_sum_0[3] ));
    XNOR3 
        \un2_d7_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_21), .B(ADD_5x5_slow_I4_Y_0_16), .C(
        \mult1_un96_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_20));
    AX1D \un2_d7_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_16), .B(ADD_5x5_slow_I3_CO1_0_15), .C(
        ADD_5x5_slow_I4_Y_2_6), .Y(\mult1_un152_sum[4] ));
    XNOR3 \un2_d3_if_generate_plus.mult1_un26_sum_ADD_4x4_slow_I3_Y_2  
        (.A(N74), .B(\rd[23]_net_1 ), .C(\mult1_un19_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_2_19));
    XNOR2 \un2_d5_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_13), .B(\mult1_un61_sum_0[4] ), .Y(
        \mult1_un68_sum_1[1] ));
    AX1D \un2_d5_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_33), .B(ADD_5x5_slow_I3_CO1_0_32), .C(
        ADD_5x5_slow_I4_Y_2_25), .Y(\mult1_un89_sum_0[4] ));
    AO1D 
        \un2_d5_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I1_CO1_1  
        (.A(\mult1_un152_sum_0[4] ), .B(\rd[3]_net_1 ), .C(
        I1_un3_CO1_3), .Y(N85_1_0));
    XOR2 \un2_d7_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_9), .B(\mult1_un89_sum[4] ), .Y(
        \mult1_un96_sum_0[1] ));
    OR2 
        \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I1_CO1_1  
        (.A(I1_un3_CO1_3), .B(I1_un2_CO1_14), .Y(N74_1_0));
    XOR2 \un2_d6_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_2), .B(N83_3), .Y(
        \mult1_un145_sum_0[3] ));
    XNOR2 \un2_d7_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1), .B(\mult1_un26_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_39));
    XA1B 
        \un2_d6_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I1_un2_CO1  
        (.A(N83_0), .B(ADD_5x5_slow_I2_S_2_10), .C(\rd[14]_net_1 ), .Y(
        I1_un2_CO1_9));
    XA1B 
        \un2_d6_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_un2_CO1  
        (.A(N83_15), .B(ADD_5x5_slow_I2_S_2), .C(\rd[2]_net_1 ), .Y(
        I1_un2_CO1_11));
    XOR2 \un2_d6_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_13), .B(N83_9), .Y(
        \mult1_un68_sum_0[3] ));
    XOR3 \un2_d5_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un26_sum_0[4] ), .B(\mult1_un26_sum_0[1] ), .C(
        N85_33), .Y(\mult1_un33_sum_0[2] ));
    NOR2B 
        \un2_d3_if_generate_plus.mult1_un61_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(N74_14), .B(\mult1_un54_sum[1] ), .Y(I2_un4_CO1_3));
    XNOR2 \un2_d5_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_8), .B(\mult1_un61_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_30));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un166_sum_ADD_4x4_slow_I1_un2_CO1  
        (.A(\mult1_un159_sum[3] ), .B(\rd[2]_net_1 ), .Y(I1_un2_CO1_0));
    AX1D \un2_d5_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_29), .B(ADD_5x5_slow_I3_CO1_0_28), .C(
        ADD_5x5_slow_I4_Y_2_13), .Y(\mult1_un138_sum_0[4] ));
    DFN1C0 \rd[17]  (.D(\rd[16]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[17]_net_1 ));
    AO13 \un2_d6_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un68_sum_0[3] ), .B(\rd[15]_net_1 ), .C(
        \rd[16]_net_1 ), .Y(N83_10));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un33_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(ADD_4x4_slow_I2_un1_CO1_0_tz_2), .B(\mult1_un26_sum[3] ), 
        .Y(ADD_4x4_slow_I2_un1_CO1_0_15));
    OR2 
        \un2_d7_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(I2_un5_CO1_2), .B(I2_un1_CO1_1_10), .Y(I2_un1_CO1_21));
    AO1 
        \un2_d3_if_generate_plus.mult1_un33_sum_ADD_4x4_slow_I2_un1_CO1  
        (.A(N74_18), .B(\mult1_un26_sum[1] ), .C(
        ADD_4x4_slow_I2_un1_CO1_0_15), .Y(I2_un1_CO1_48));
    XNOR3 
        \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I3_Y_2  
        (.A(I2_un1_CO1_18), .B(ADD_4x4_slow_I3_Y_2_0), .C(
        ADD_4x4_slow_I3_Y_1_0), .Y(ADD_4x4_slow_I3_Y_2_1));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_21), .B(\mult1_un117_sum[2] ), .C(
        \mult1_un117_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_33));
    XOR3 \un2_d5_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un152_sum_0[4] ), .B(\mult1_un152_sum_1[1] ), .C(
        N85_36), .Y(\mult1_un159_sum_0[2] ));
    XOR2 \un2_d7_if_generate_plus.mult1_un1_sum_I_7  (.A(
        ADD_5x5_slow_I1_S_1), .B(ADD_5x5_slow_I4_Y_0_27), .Y(
        \DWACT_ADD_CI_0_pog_array_0[0] ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(\mult1_un166_sum[1] ), .B(N85_35), .Y(I2_un4_CO1_15));
    XOR2 \un2_d6_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_15), .B(\mult1_un54_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_13));
    DFN1E1 \cur_rand_1[3]  (.D(\d2[0]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[3]));
    AO13 \un2_d7_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un33_sum[4] ), .B(\rd[19]_net_1 ), .C(
        \rd[20]_net_1 ), .Y(N85_14));
    AO1 
        \un2_d3_if_generate_plus.mult1_un26_sum_ADD_4x4_slow_I2_un1_CO1  
        (.A(N74_19), .B(\mult1_un19_sum_0[1] ), .C(
        ADD_4x4_slow_I2_un1_CO1_0_16), .Y(I2_un1_CO1_47));
    AO13 
        \un2_d3_if_generate_plus.mult1_un117_sum_ADD_4x4_slow_I2_un1_CO1  
        (.A(N74_6), .B(\mult1_un110_sum_0[1] ), .C(
        \mult1_un110_sum[3] ), .Y(I2_un1_CO1_42));
    XNOR2 
        \un2_d5_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un89_sum_0[2] ), .B(\mult1_un89_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_18));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(\mult1_un159_sum[1] ), .B(N85_18), .Y(I2_un4_CO1_14));
    XOR2 \un2_d6_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_16), .B(\mult1_un47_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_14));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un26_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(I1_un3_CO1_13), .B(\mult1_un19_sum_0[1] ), .C(
        \mult1_un19_sum[3] ), .Y(ADD_4x4_slow_I2_un1_CO1_0_16));
    AX1D \un2_d3_if_generate_plus.mult1_un89_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_1), .B(ADD_4x4_slow_I2_un1_CO1_0), .C(
        ADD_4x4_slow_I3_Y_2_10), .Y(\mult1_un89_sum[3] ));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un40_sum_ADD_4x4_slow_I1_CO1_1  
        (.A(\rd[19]_net_1 ), .B(\mult1_un33_sum[3] ), .C(
        \rd[20]_net_1 ), .Y(N74_1_9));
    XOR2 \un2_d7_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_3), .B(\mult1_un131_sum[4] ), .Y(
        \mult1_un138_sum[1] ));
    XOR2 \un2_d3_if_generate_plus.mult1_un33_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_18), .B(\mult1_un26_sum[3] ), .Y(
        \mult1_un33_sum[1] ));
    XOR3 \un2_d7_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un47_sum[4] ), .B(\mult1_un47_sum_0[1] ), .C(N85_13), 
        .Y(\mult1_un54_sum[2] ));
    XOR2 \un2_d7_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_6), .B(\mult1_un110_sum[4] ), .Y(
        \mult1_un117_sum_1[1] ));
    OR2 
        \un2_d5_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(I2_un5_CO1_4), .B(I2_un1_CO1_1_13), .Y(I2_un1_CO1_33));
    XA1A 
        \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(I2_un1_CO1_18), .B(ADD_4x4_slow_I3_Y_2_0), .C(
        ADD_4x4_slow_I2_un1_CO1_0_tz), .Y(ADD_4x4_slow_I2_un1_CO1_0_4));
    AX1D \un2_d7_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_5), .B(ADD_5x5_slow_I3_CO1_0_4), .C(
        ADD_5x5_slow_I4_Y_2_37), .Y(\mult1_un40_sum[4] ));
    NOR2 \d6_RNO[2]  (.A(reset_c), .B(I_14_4), .Y(\d6_RNO[2]_net_1 ));
    XNOR3 
        \un2_d3_if_generate_plus.mult1_un110_sum_ADD_4x4_slow_I3_Y_1  
        (.A(\mult1_un96_sum[3] ), .B(\mult1_un96_sum[1] ), .C(N74_8), 
        .Y(ADD_4x4_slow_I3_Y_1_5));
    XOR2 \un2_d7_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_0_6), .B(N85_26), .Y(\mult1_un117_sum[2] )
        );
    XOR3 \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I2_S_0  
        (.A(\mult1_un159_sum[4] ), .B(ADD_4x4_slow_I1_S_0), .C(
        \mult1_un166_sum[4] ), .Y(ADD_5x5_slow_I2_S_0));
    XOR3 \un2_d7_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un124_sum[4] ), .B(\mult1_un124_sum_1[1] ), .C(
        N85_22), .Y(\mult1_un131_sum[2] ));
    XNOR2 \un2_d5_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I1_S  
        (.A(ADD_4x4_slow_I1_S_0), .B(\mult1_un159_sum_0[4] ), .Y(
        \mult1_un166_sum[1] ));
    XNOR2 
        \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un131_sum_0[2] ), .B(\mult1_un131_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_9));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(\mult1_un117_sum_1[1] ), .B(N85_24), .Y(I2_un4_CO1_21));
    DFN1C0 \rd[18]  (.D(\rd[17]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[18]_net_1 ));
    XOR3 \un2_d6_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I1_S  (
        .A(N83), .B(ADD_5x5_slow_I2_S_2_0), .C(ADD_4x4_slow_I1_S_0_1), 
        .Y(\mult1_un166_sum_0[2] ));
    XOR2 \un2_d6_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_7), .B(\mult1_un110_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_5));
    XOR2 \un2_d7_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_17), .B(\mult1_un33_sum[4] ), .Y(
        \mult1_un40_sum_0[1] ));
    OA1 
        \un2_d7_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(N85_15), .B(\mult1_un131_sum[4] ), .C(
        \mult1_un131_sum_0[1] ), .Y(I2_un1_CO1_1_5));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_17), .B(\mult1_un103_sum[2] ), .Y(I3_un3_CO1_21)
        );
    XOR2 \un2_d3_if_generate_plus.mult1_un47_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_16), .B(\mult1_un40_sum[3] ), .Y(
        \mult1_un47_sum[1] ));
    XNOR2 
        \un2_d6_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_5), .B(\mult1_un117_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_5));
    AO1 \un2_d3_if_generate_plus.mult1_un40_sum_ADD_4x4_slow_I1_CO1  (
        .A(\mult1_un33_sum[3] ), .B(\rd[19]_net_1 ), .C(N74_1_9), .Y(
        N74_17));
    NOR2A \un2_d7_if_generate_plus.mult1_un1_sum_I_1  (.A(
        ADD_5x5_slow_I4_Y_0_27), .B(\rd[0]_net_1 ), .Y(
        \DWACT_ADD_CI_0_TMP_0[0] ));
    XNOR2 \un2_d5_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_18), .B(\mult1_un26_sum_0[4] ), .Y(
        \mult1_un33_sum_1[1] ));
    NOR2A \un2_d5_if_generate_plus.mult1_un19_sum_ADD_5x5_slow_I1_CO1  
        (.A(\rd[22]_net_1 ), .B(\rd[23]_net_1 ), .Y(N85_1));
    AO1 \un2_d3_if_generate_plus.mult1_un75_sum_ADD_4x4_slow_I1_CO1  (
        .A(\mult1_un68_sum[3] ), .B(\rd[14]_net_1 ), .C(N74_1_5), .Y(
        N74_12));
    OR2 
        \un2_d5_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(ADD_5x5_slow_I2_un1_CO1_0_14), .B(I2_un4_CO1_31), .Y(
        I2_un1_CO1_40));
    AX1D \un2_d3_if_generate_plus.mult1_un61_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_3), .B(ADD_4x4_slow_I2_un1_CO1_0_1), .C(
        ADD_4x4_slow_I3_Y_2_14), .Y(\mult1_un61_sum[3] ));
    OR2 
        \un2_d5_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(ADD_5x5_slow_I2_un1_CO1_0_1), .B(I2_un4_CO1_18), .Y(
        I2_un1_CO1_6));
    XNOR2 \un2_d5_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I1_S  
        (.A(ADD_4x4_slow_I1_S_0_3), .B(\mult1_un131_sum_0[4] ), .Y(
        \mult1_un138_sum_0[1] ));
    XNOR3 \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_28), .B(ADD_5x5_slow_I4_Y_0_21), .C(
        \mult1_un75_sum_0[4] ), .Y(ADD_5x5_slow_I4_Y_2_26));
    NOR2A \d6_RNO_0[2]  (.A(I_14_4), .B(reset_c), .Y(
        \d6_RNO_0[2]_net_1 ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(\mult1_un61_sum_0[4] ), .B(ADD_5x5_slow_I2_un1_CO1_0_tz_1), 
        .Y(ADD_5x5_slow_I2_un1_CO1_0_9));
    XNOR2 \un2_d6_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_14), .B(\mult1_un54_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_14));
    XA1A 
        \un2_d6_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(N83_15), .B(ADD_5x5_slow_I2_S_2), .C(
        ADD_5x5_slow_I2_un1_CO1_0_tz_0), .Y(
        ADD_5x5_slow_I2_un1_CO1_0_8));
    NOR2B 
        \un2_d3_if_generate_plus.mult1_un145_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(N74_2), .B(\mult1_un138_sum_1[1] ), .Y(I2_un4_CO1_5));
    MAJ3 
        \un2_d7_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\mult1_un47_sum_0[1] ), .B(\mult1_un47_sum[4] ), .C(N85_13)
        , .Y(I2_un1_CO1_32));
    XNOR3 
        \un2_d7_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_3), .B(ADD_5x5_slow_I4_Y_0_0), .C(
        \mult1_un159_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_2));
    XNOR2 \un2_d3_if_generate_plus.mult1_un54_sum_ADD_4x4_slow_I3_Y_0  
        (.A(\mult1_un40_sum[1] ), .B(\mult1_un40_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_0_10));
    XNOR3 
        \un2_d3_if_generate_plus.mult1_un131_sum_ADD_4x4_slow_I3_Y_1  
        (.A(\mult1_un117_sum[3] ), .B(\mult1_un117_sum[1] ), .C(N74_5), 
        .Y(ADD_4x4_slow_I3_Y_1_2));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un138_sum_ADD_4x4_slow_I3_Y_2  
        (.A(ADD_4x4_slow_I3_Y_1_1), .B(\mult1_un131_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_2_3));
    XNOR2 
        \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_3), .B(\mult1_un117_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_17));
    MAJ3 
        \un2_d7_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\mult1_un138_sum[4] ), .B(N85_23), .C(\mult1_un138_sum[1] )
        , .Y(I2_un1_CO1_7));
    XOR3 \un2_d5_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un124_sum_0[4] ), .B(\mult1_un124_sum_0[1] ), .C(
        N85_16), .Y(\mult1_un131_sum_0[2] ));
    AX1D \un2_d7_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_4), .B(ADD_5x5_slow_I3_CO1_0_3), .C(
        ADD_5x5_slow_I4_Y_2_27), .Y(\mult1_un75_sum_0[4] ));
    NOR2A \d3_RNO_0[0]  (.A(\DWACT_ADD_CI_0_partial_sum_1[0] ), .B(
        reset_c), .Y(\d3_RNO_0[0]_net_1 ));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_15), .B(\mult1_un26_sum[2] ), .C(
        \mult1_un26_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_36));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_24), .B(\mult1_un89_sum_0[2] ), .C(
        \mult1_un89_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_31));
    DFN1E1 \cur_rand_1[14]  (.D(\d5[2]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[14]));
    XOR2 \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I4_Y  (
        .A(ADD_5x5_slow_I4_Y_2_26), .B(N89_1), .Y(
        \mult1_un82_sum_0[4] ));
    XOR2 \un2_d7_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_16), .B(\mult1_un40_sum[4] ), .Y(
        \mult1_un47_sum_0[1] ));
    AO13 \un2_d6_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un89_sum_0[3] ), .B(\rd[12]_net_1 ), .C(
        \rd[13]_net_1 ), .Y(N83_18));
    XNOR3 
        \un2_d7_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_7), .B(ADD_5x5_slow_I4_Y_0_4), .C(
        \mult1_un145_sum_0[4] ), .Y(ADD_5x5_slow_I4_Y_2_6));
    XOR2 \un2_d6_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_4), .B(N83_5), .Y(
        \mult1_un131_sum_0[3] ));
    NOR2 \d4_RNO[1]  (.A(reset_c), .B(\rd[1]_net_1 ), .Y(
        \d4_RNO[1]_net_1 ));
    XNOR2 
        \un2_d6_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_7), .B(\mult1_un103_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_7));
    XNOR2 \un2_d5_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un47_sum_0[2] ), .B(\mult1_un47_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_25));
    AX1D \un2_d5_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I4_Y_1  
        (.A(I2_un1_CO1_1_2), .B(I2_un5_CO1_1), .C(
        ADD_5x5_slow_I4_Y_0_24), .Y(ADD_5x5_slow_I4_Y_1_8));
    NOR2A 
        \un2_d5_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(ADD_5x5_slow_I3_CO1_0_tz_0), .B(\mult1_un96_sum_0[4] ), .Y(
        ADD_5x5_slow_I3_CO1_0_34));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un47_sum_ADD_4x4_slow_I1_CO1_1  
        (.A(\mult1_un40_sum[3] ), .B(\rd[18]_net_1 ), .C(
        \rd[19]_net_1 ), .Y(N74_1_8));
    NOR2A 
        \un2_d5_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I1_un3_CO1  
        (.A(\rd[14]_net_1 ), .B(\rd[15]_net_1 ), .Y(I1_un3_CO1_14));
    AO1 \un2_d3_if_generate_plus.mult1_un138_sum_ADD_4x4_slow_I1_CO1  
        (.A(\mult1_un131_sum[3] ), .B(\rd[5]_net_1 ), .C(N74_1_1), .Y(
        N74_3));
    XNOR2 \un2_d3_if_generate_plus.mult1_un68_sum_ADD_4x4_slow_I3_Y_0  
        (.A(\mult1_un54_sum[1] ), .B(\mult1_un54_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_0_8));
    XOR2 \un2_d6_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_12), .B(\mult1_un75_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_10));
    AO13 \un2_d3_if_generate_plus.mult1_un96_sum_ADD_4x4_slow_I1_CO1  
        (.A(\mult1_un89_sum[3] ), .B(\rd[11]_net_1 ), .C(
        \rd[12]_net_1 ), .Y(N74_9));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_39), .B(\mult1_un26_sum_0[2] ), .Y(
        I3_un3_CO1_26));
    OR2 \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I3_CO1  (
        .A(I3_un3_CO1_1), .B(ADD_5x5_slow_I3_CO1_0_0), .Y(N89));
    XNOR2 \un2_d5_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_15), .B(\mult1_un26_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_40));
    XNOR3 
        \un2_d3_if_generate_plus.mult1_un103_sum_ADD_4x4_slow_I3_Y_1  
        (.A(\mult1_un89_sum[3] ), .B(\mult1_un89_sum[1] ), .C(N74_9), 
        .Y(ADD_4x4_slow_I3_Y_1_6));
    XNOR2 \un2_d5_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I1_S  
        (.A(ADD_4x4_slow_I1_S_0_6), .B(\mult1_un110_sum_0[4] ), .Y(
        \mult1_un117_sum_0[1] ));
    AX1D \un2_d5_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_25), .B(ADD_5x5_slow_I3_CO1_0_24), .C(
        ADD_5x5_slow_I4_Y_2_28), .Y(\mult1_un75_sum[4] ));
    AX1D \un2_d7_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_18), .B(ADD_5x5_slow_I3_CO1_0_17), .C(
        ADD_5x5_slow_I4_Y_2_8), .Y(\mult1_un145_sum_0[4] ));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_31), .B(\mult1_un19_sum_0[2] ), .C(
        \mult1_un19_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_26));
    XOR3 \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_S  (
        .A(\rd[1]_net_1 ), .B(\rd[0]_net_1 ), .C(
        \mult1_un166_sum_0[4] ), .Y(ADD_5x5_slow_I1_S));
    OA1 
        \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_1_3), .B(I2_un5_CO1_3), .C(\mult1_un166_sum[2] )
        , .Y(I3_un3_CO1_13));
    XNOR3 \un2_d3_if_generate_plus.mult1_un68_sum_ADD_4x4_slow_I3_Y_2  
        (.A(N74_14), .B(ADD_4x4_slow_I3_Y_0_8), .C(\mult1_un61_sum[3] )
        , .Y(ADD_4x4_slow_I3_Y_2_13));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un103_sum_ADD_4x4_slow_I3_Y_2  
        (.A(ADD_4x4_slow_I3_Y_1_6), .B(\mult1_un96_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_2_8));
    AO13 \un2_d7_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un47_sum[4] ), .B(\rd[17]_net_1 ), .C(
        \rd[18]_net_1 ), .Y(N85_13));
    XNOR2 \un2_d3_if_generate_plus.mult1_un82_sum_ADD_4x4_slow_I3_Y_0  
        (.A(\mult1_un68_sum[1] ), .B(\mult1_un68_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_0_7));
    XOR3 \un2_d5_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un110_sum_0[4] ), .B(\mult1_un110_sum_1[1] ), .C(
        N85_27), .Y(\mult1_un117_sum_0[2] ));
    NOR2B 
        \un2_d3_if_generate_plus.mult1_un89_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(N74_10), .B(\mult1_un82_sum_0[1] ), .Y(I2_un4_CO1_1));
    XOR2 \un2_d6_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_6), .B(N83_7), .Y(
        \mult1_un117_sum_0[3] ));
    XNOR3 
        \un2_d5_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_8), .B(ADD_5x5_slow_I4_Y_0_5), .C(
        \mult1_un152_sum_0[4] ), .Y(ADD_5x5_slow_I4_Y_2_7));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un40_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(N74_1_9), .B(\mult1_un33_sum[1] ), .C(\mult1_un33_sum[3] ), 
        .Y(ADD_4x4_slow_I2_un1_CO1_0_9));
    XNOR3 
        \un2_d3_if_generate_plus.mult1_un166_sum_ADD_4x4_slow_I3_Y_0  
        (.A(I2_un1_CO1_18), .B(ADD_4x4_slow_I3_Y_2_0), .C(
        \mult1_un152_sum_0[1] ), .Y(ADD_4x4_slow_I3_Y_0_0));
    DFN1P1C1 \d2[0]  (.D(\rd[0]_net_1 ), .CLK(ref_signal_c), .PRE(
        \d2_RNO_0[0]_net_1 ), .CLR(\d2_RNO[0]_net_1 ), .Q(
        \d2[0]_net_1 ));
    XNOR2 
        \un2_d7_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un110_sum[2] ), .B(\mult1_un110_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_12));
    AO13 \un2_d7_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I3_CO1  
        (.A(I2_un1_CO1_19), .B(\mult1_un96_sum[2] ), .C(
        \mult1_un96_sum[4] ), .Y(N89_6));
    AO1 
        \un2_d5_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N85_32), .B(\mult1_un61_sum_1[1] ), .C(
        ADD_5x5_slow_I2_un1_CO1_0_9), .Y(I2_un1_CO1_30));
    AXOI5 
        \un2_d6_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(\rd[21]_net_1 ), .B(\rd[22]_net_1 ), .C(\rd[23]_net_1 ), 
        .Y(I2_un4_CO1_0));
    AO1D 
        \un2_d5_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I1_CO1_1  
        (.A(\mult1_un82_sum[4] ), .B(\rd[13]_net_1 ), .C(I1_un3_CO1_0), 
        .Y(N85_1_2));
    AX1D \un2_d7_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_2), .B(ADD_5x5_slow_I3_CO1_0_1), .C(
        ADD_5x5_slow_I4_Y_2_22), .Y(\mult1_un96_sum[4] ));
    XNOR2 
        \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un159_sum[2] ), .B(\mult1_un159_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0));
    AO14 \un2_d6_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I2_S_3  
        (.A(\rd[22]_net_1 ), .B(\rd[21]_net_1 ), .C(\rd[23]_net_1 ), 
        .Y(ADD_5x5_slow_I2_S_3));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un117_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[8]_net_1 ), .B(\rd[9]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_6));
    AX1D \un2_d7_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_6), .B(ADD_5x5_slow_I3_CO1_0_5), .C(
        ADD_5x5_slow_I4_Y_2_35), .Y(\mult1_un47_sum[4] ));
    DFN1C0 \rd[15]  (.D(\rd[14]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[15]_net_1 ));
    XNOR3 \un2_d5_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_27), .B(ADD_5x5_slow_I4_Y_0_20), .C(
        \mult1_un82_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_25));
    XOR3 \un2_d7_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un61_sum[4] ), .B(\mult1_un61_sum_0[1] ), .C(N85_6), 
        .Y(\mult1_un68_sum[2] ));
    AO18 \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un138_sum_0[4] ), .B(\rd[4]_net_1 ), .C(
        \rd[5]_net_1 ), .Y(N85_37));
    AO13 \un2_d3_if_generate_plus.mult1_un117_sum_ADD_4x4_slow_I1_CO1  
        (.A(\mult1_un110_sum[3] ), .B(\rd[8]_net_1 ), .C(\rd[9]_net_1 )
        , .Y(N74_6));
    AO1 \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I3_CO1  (
        .A(I2_un1_CO1_26), .B(\mult1_un75_sum[2] ), .C(
        ADD_5x5_slow_I3_CO1_0_35), .Y(N89_1));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_38), .B(\mult1_un26_sum[2] ), .Y(I3_un3_CO1_36));
    XOR2 \un2_d7_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I2_S_0  
        (.A(\mult1_un103_sum[1] ), .B(\mult1_un103_sum[4] ), .Y(
        ADD_5x5_slow_I2_S_0_7));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_13), .B(\mult1_un47_sum_0[2] ), .C(
        \mult1_un47_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_21));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un138_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(N74_1_1), .B(\mult1_un131_sum[1] ), .C(
        \mult1_un131_sum[3] ), .Y(ADD_4x4_slow_I2_un1_CO1_0_2));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_2), .B(\mult1_un159_sum[2] ), .Y(I3_un3_CO1_12));
    XOR2 \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_0_5), .B(N85_37), .Y(
        \mult1_un145_sum_0[2] ));
    XOR2 \un2_d7_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I4_Y  (
        .A(I2_un1_CO1), .B(I3_un3_CO1), .Y(\mult1_un26_sum[4] ));
    XNOR2 \un2_d7_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_7), .B(\mult1_un61_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_29));
    XNOR2 
        \un2_d6_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_1), .B(\mult1_un145_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_1));
    XOR3 \un2_d5_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un61_sum_0[4] ), .B(\mult1_un61_sum_1[1] ), .C(
        N85_32), .Y(\mult1_un68_sum_0[2] ));
    DFN1E1 \cur_rand_1[6]  (.D(\d3[0]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[6]));
    XNOR2 \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_1), .B(\mult1_un82_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_0));
    NOR2B 
        \un2_d3_if_generate_plus.mult1_un110_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(N74_7), .B(\mult1_un103_sum_0[1] ), .Y(I2_un4_CO1_10));
    XOR2 \un2_d3_if_generate_plus.mult1_un40_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_17), .B(\mult1_un33_sum[3] ), .Y(
        \mult1_un40_sum[1] ));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_0), .B(\mult1_un19_sum[2] ), .Y(I3_un3_CO1));
    AO1 
        \un2_d5_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I3_CO1_0_tz  
        (.A(N85_39), .B(\mult1_un96_sum_1[1] ), .C(
        \mult1_un96_sum_0[2] ), .Y(ADD_5x5_slow_I3_CO1_0_tz_0));
    XOR2 \un2_d3_if_generate_plus.mult1_un124_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_5), .B(\mult1_un117_sum[3] ), .Y(
        \mult1_un124_sum[1] ));
    XNOR2 \un2_d3_if_generate_plus.mult1_un96_sum_ADD_4x4_slow_I3_Y_0  
        (.A(\mult1_un82_sum_0[1] ), .B(\mult1_un82_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_0_5));
    AX1D \un2_d3_if_generate_plus.mult1_un47_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_12), .B(ADD_4x4_slow_I2_un1_CO1_0_10), .C(
        ADD_4x4_slow_I3_Y_2_16), .Y(\mult1_un47_sum[3] ));
    XNOR2 \un2_d3_if_generate_plus.mult1_un75_sum_ADD_4x4_slow_I3_Y_2  
        (.A(ADD_4x4_slow_I3_Y_1_7), .B(\mult1_un68_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_2_12));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un145_sum_ADD_4x4_slow_I1_un2_CO1  
        (.A(\mult1_un138_sum[3] ), .B(\rd[5]_net_1 ), .Y(I1_un2_CO1_5));
    NOR2A \d6_RNO_0[1]  (.A(\DWACT_ADD_CI_0_partial_sum[1] ), .B(
        reset_c), .Y(\d6_RNO_0[1]_net_1 ));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_6), .B(\mult1_un124_sum[2] ), .C(
        \mult1_un124_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_6));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_3), .B(\mult1_un166_sum[2] ), .C(
        \mult1_un166_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_12));
    MAJ3 
        \un2_d7_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\mult1_un96_sum_0[1] ), .B(\mult1_un96_sum[4] ), .C(N85_9), 
        .Y(I2_un1_CO1_19));
    OA1 
        \un2_d5_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(I1_un3_CO1_9), .B(\mult1_un89_sum_1[1] ), .C(
        \mult1_un89_sum_0[4] ), .Y(ADD_5x5_slow_I2_un1_CO1_0_6));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un145_sum_ADD_4x4_slow_I3_Y_0  
        (.A(\mult1_un131_sum[1] ), .B(\mult1_un131_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_0_3));
    AO1 
        \un2_d7_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N85_22), .B(\mult1_un124_sum[4] ), .C(I2_un1_CO1_1_6), .Y(
        I2_un1_CO1_11));
    NOR2A \d5_RNO_0[1]  (.A(I_12_4), .B(reset_c), .Y(
        \d5_RNO_0[1]_net_1 ));
    XNOR3 \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_S  
        (.A(\rd[1]_net_1 ), .B(\rd[0]_net_1 ), .C(\mult1_un166_sum[4] )
        , .Y(ADD_5x5_slow_I1_S_1));
    AO13 \un2_d6_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un103_sum_0[3] ), .B(\rd[10]_net_1 ), .C(
        \rd[11]_net_1 ), .Y(N83_16));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(N85_41), .B(\mult1_un89_sum_1[1] ), .Y(I2_un4_CO1_24));
    NOR2A 
        \un2_d5_if_generate_plus.mult1_un19_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(N85_1), .B(\rd[23]_net_1 ), .Y(I2_un4_CO1));
    XOR2 \un2_d3_if_generate_plus.mult1_un103_sum_ADD_4x4_slow_I3_Y  (
        .A(ADD_4x4_slow_I3_Y_2_8), .B(I2_un1_CO1_45), .Y(
        \mult1_un103_sum[3] ));
    DFN1C0 \rd[21]  (.D(\rd[20]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[21]_net_1 ));
    DFN1C0 \rd[12]  (.D(\rd[11]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[12]_net_1 ));
    NOR2 
        \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I1_un2_CO1  
        (.A(\mult1_un145_sum[4] ), .B(\rd[4]_net_1 ), .Y(I1_un2_CO1));
    AO18 \un2_d5_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un103_sum_0[4] ), .B(\rd[9]_net_1 ), .C(
        \rd[10]_net_1 ), .Y(N85_40));
    OR2 \un2_d3_if_generate_plus.mult1_un82_sum_ADD_4x4_slow_I1_CO1  (
        .A(ADD_4x4_slow_I1_CO1_0_2), .B(I1_un2_CO1_3), .Y(N74_11));
    XNOR2 \un2_d3_if_generate_plus.mult1_un47_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[18]_net_1 ), .B(\rd[19]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_16));
    XOR2 \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_0_8), .B(N85_4), .Y(\mult1_un89_sum[2] ));
    XOR2 \un2_d7_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_2), .B(\mult1_un145_sum_0[4] ), .Y(
        \mult1_un152_sum[1] ));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_12), .B(\mult1_un75_sum_0[2] ), .C(
        \mult1_un75_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0));
    AO1 \un2_d3_if_generate_plus.mult1_un124_sum_ADD_4x4_slow_I1_CO1  
        (.A(\mult1_un117_sum[3] ), .B(\rd[7]_net_1 ), .C(N74_1_2), .Y(
        N74_5));
    AO18 \un2_d5_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un19_sum[4] ), .B(\rd[21]_net_1 ), .C(
        \rd[22]_net_1 ), .Y(N85_12));
    XOR2 \un2_d7_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_8), .B(\mult1_un96_sum[4] ), .Y(
        \mult1_un103_sum[1] ));
    XOR2 \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I2_S_0  
        (.A(\mult1_un138_sum_0[1] ), .B(\mult1_un138_sum_0[4] ), .Y(
        ADD_5x5_slow_I2_S_0_5));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I2_un5_CO1  
        (.A(I1_un3_CO1_1), .B(\mult1_un75_sum[4] ), .Y(I2_un5_CO1_5));
    XOR3 \un2_d5_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un54_sum_0[4] ), .B(\mult1_un54_sum_1[1] ), .C(
        N85_29), .Y(\mult1_un61_sum_0[2] ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(\mult1_un131_sum_1[1] ), .B(I2_un1_CO1_1_tz_4), .Y(
        I2_un1_CO1_1_7));
    XOR2 \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I2_S_0  
        (.A(\mult1_un75_sum[1] ), .B(\mult1_un75_sum_0[4] ), .Y(
        ADD_5x5_slow_I2_S_0_9));
    OR3 \un2_d6_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I1_CO1  (
        .A(I1_un5_CO1_0), .B(I1_un3_CO1_1), .C(I1_un2_CO1_9), .Y(
        N83_12));
    NOR3B 
        \un2_d5_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I2_un5_CO1  
        (.A(\rd[17]_net_1 ), .B(\mult1_un47_sum_0[4] ), .C(
        \rd[18]_net_1 ), .Y(I2_un5_CO1_4));
    AO13 \un2_d7_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un145_sum_0[4] ), .B(\rd[3]_net_1 ), .C(
        \rd[4]_net_1 ), .Y(N85_19));
    AO13 \un2_d3_if_generate_plus.mult1_un173_sum_ADD_4x4_slow_I1_CO1  
        (.A(\mult1_un166_sum[3] ), .B(\rd[0]_net_1 ), .C(\rd[1]_net_1 )
        , .Y(N74_20));
    XNOR2 
        \un2_d5_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un103_sum_0[2] ), .B(\mult1_un103_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_15));
    AND2 
        \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(I2_un1_CO1_1_tz), .B(\mult1_un145_sum[1] ), .Y(
        I2_un1_CO1_1));
    AX1D \un2_d7_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_19), .B(ADD_5x5_slow_I3_CO1_0_18), .C(
        ADD_5x5_slow_I4_Y_2_16), .Y(\mult1_un117_sum[4] ));
    AOI1 
        \un2_d6_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N83_14), .B(\mult1_un166_sum_0[2] ), .C(
        ADD_5x5_slow_I2_un1_CO1_0_8), .Y(I2_un1_CO1_49));
    XNOR3 \un2_d3_if_generate_plus.mult1_un173_sum_ADD_4x4_slow_I1_S  
        (.A(\rd[1]_net_1 ), .B(\rd[0]_net_1 ), .C(\mult1_un166_sum[3] )
        , .Y(ADD_4x4_slow_I1_S));
    DFN1P1C1 \d8[2]  (.D(\rd[2]_net_1 ), .CLK(ref_signal_c), .PRE(
        \d8_RNO_0[2]_net_1 ), .CLR(\d8_RNO[2]_net_1 ), .Q(
        \d8[2]_net_1 ));
    AO13 \un2_d7_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un110_sum[4] ), .B(\rd[8]_net_1 ), .C(\rd[9]_net_1 )
        , .Y(N85_26));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_24), .B(\mult1_un89_sum_0[2] ), .Y(
        I3_un3_CO1_32));
    XNOR2 \un2_d6_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_12), .B(\mult1_un68_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_2_12));
    NOR2A 
        \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I1_un2_CO1  
        (.A(\mult1_un75_sum_0[4] ), .B(\rd[14]_net_1 ), .Y(
        I1_un2_CO1_1));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1), .B(\mult1_un145_sum_0[2] ), .C(
        \mult1_un145_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_27));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un26_sum_ADD_4x4_slow_I1_un3_CO1  
        (.A(\rd[21]_net_1 ), .B(\rd[22]_net_1 ), .Y(I1_un3_CO1_13));
    DFN1C0 \rd[23]  (.D(\rd[22]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[23]_net_1 ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(\mult1_un159_sum_1[1] ), .B(N85_20), .Y(I2_un4_CO1_16));
    AO1A \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un117_sum_0[4] ), .B(\rd[7]_net_1 ), .C(N85_1_1), 
        .Y(N85_17));
    AX1D \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_11), .B(ADD_5x5_slow_I3_CO1_0_10), .C(
        ADD_5x5_slow_I4_Y_2_4), .Y(\mult1_un159_sum[4] ));
    AO13 \un2_d7_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un117_sum[4] ), .B(\rd[7]_net_1 ), .C(\rd[8]_net_1 )
        , .Y(N85_24));
    AX1D \un2_d3_if_generate_plus.mult1_un124_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_9), .B(ADD_4x4_slow_I2_un1_CO1_0_7), .C(
        ADD_4x4_slow_I3_Y_2_5), .Y(\mult1_un124_sum[3] ));
    XNOR2 \un2_d3_if_generate_plus.mult1_un89_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[12]_net_1 ), .B(\rd[13]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_10));
    AX1D \un2_d5_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_26), .B(ADD_5x5_slow_I3_CO1_0_25), .C(
        ADD_5x5_slow_I4_Y_2_40), .Y(\mult1_un33_sum_0[4] ));
    NOR2A \un2_d5_if_generate_plus.mult1_un1_sum_I_1  (.A(
        ADD_5x5_slow_I4_Y), .B(\rd[0]_net_1 ), .Y(
        \DWACT_ADD_CI_0_TMP[0] ));
    XNOR2 
        \un2_d7_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un89_sum[2] ), .B(\mult1_un89_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_16));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_1), .B(\mult1_un68_sum_0[2] ), .C(
        \mult1_un68_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_24));
    XOR3 \un2_d7_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un145_sum_0[4] ), .B(\mult1_un145_sum_0[1] ), .C(
        N85_19), .Y(\mult1_un152_sum[2] ));
    XNOR3 
        \un2_d5_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_6), .B(ADD_5x5_slow_I4_Y_0_3), .C(
        \mult1_un159_sum_0[4] ), .Y(ADD_5x5_slow_I4_Y_2_5));
    NOR2 \d3_RNO[1]  (.A(reset_c), .B(I_10), .Y(\d3_RNO[1]_net_1 ));
    XNOR2 \rd_RNO[0]  (.A(\rd[23]_net_1 ), .B(\rd[11]_net_1 ), .Y(
        \rd_RNO[0]_net_1 ));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un117_sum_ADD_4x4_slow_I3_Y_2  
        (.A(ADD_4x4_slow_I3_Y_1_4), .B(\mult1_un110_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_2_6));
    XNOR3 \un2_d5_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un19_sum[4] ), .B(\mult1_un19_sum_0[2] ), .C(
        I2_un1_CO1_40), .Y(ADD_5x5_slow_I4_Y_1_15));
    AO13 \un2_d7_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un96_sum[4] ), .B(\rd[10]_net_1 ), .C(
        \rd[11]_net_1 ), .Y(N85_9));
    AX1D \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_10), .B(ADD_5x5_slow_I3_CO1_0_9), .C(
        ADD_5x5_slow_I4_Y_2_17), .Y(\mult1_un124_sum_0[4] ));
    OA1 
        \un2_d5_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_1_1), .B(I2_un5_CO1_0), .C(
        \mult1_un68_sum_0[2] ), .Y(I3_un3_CO1_25));
    AO13 \un2_d6_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un96_sum_0[3] ), .B(\rd[11]_net_1 ), .C(
        \rd[12]_net_1 ), .Y(N83_17));
    NOR2B 
        \un2_d3_if_generate_plus.mult1_un124_sum_ADD_4x4_slow_I2_un4_CO1  
        (.A(N74_5), .B(\mult1_un117_sum[1] ), .Y(I2_un4_CO1_9));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(\mult1_un61_sum_0[1] ), .B(N85_6), .Y(I2_un4_CO1_27));
    NOR2A \d3_RNO_0[1]  (.A(I_10), .B(reset_c), .Y(\d3_RNO_0[1]_net_1 )
        );
    XOR2 \un2_d7_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_14), .B(\mult1_un54_sum[4] ), .Y(
        \mult1_un61_sum_0[1] ));
    XOR2 \un2_d3_if_generate_plus.mult1_un1_sum_I_10  (.A(
        \DWACT_ADD_CI_0_partial_sum_1[1] ), .B(
        \DWACT_ADD_CI_0_TMP_1[0] ), .Y(I_10));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_16), .B(\mult1_un159_sum_0[2] ), .C(
        \mult1_un159_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_29));
    AO18 \un2_d5_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un47_sum_0[4] ), .B(\rd[17]_net_1 ), .C(
        \rd[18]_net_1 ), .Y(N85_31));
    OR2 
        \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(I2_un5_CO1_6), .B(I2_un1_CO1_1), .Y(I2_un1_CO1_8));
    XNOR2 \un2_d5_if_generate_plus.mult1_un103_sum_ADD_5x5_slow_I1_S  
        (.A(ADD_4x4_slow_I1_S_0_8), .B(\mult1_un96_sum_0[4] ), .Y(
        \mult1_un103_sum_1[1] ));
    XNOR2 \un2_d3_if_generate_plus.mult1_un61_sum_ADD_4x4_slow_I3_Y_0  
        (.A(\mult1_un47_sum[1] ), .B(\mult1_un47_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_0_9));
    XOR2 \un2_d3_if_generate_plus.mult1_un117_sum_ADD_4x4_slow_I3_Y  (
        .A(ADD_4x4_slow_I3_Y_2_6), .B(I2_un1_CO1_42), .Y(
        \mult1_un117_sum[3] ));
    OA1 
        \un2_d5_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_1_2), .B(I2_un5_CO1_1), .C(
        \mult1_un54_sum_0[2] ), .Y(I3_un3_CO1_24));
    NOR2A \d4_RNO_0[1]  (.A(\rd[1]_net_1 ), .B(reset_c), .Y(
        \d4_RNO_0[1]_net_1 ));
    XNOR2 \un2_d5_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_13), .B(\mult1_un40_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_36));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un124_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[7]_net_1 ), .B(\rd[8]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_5));
    XOR2 \un2_d7_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_0), .B(\mult1_un138_sum[4] ), .Y(
        \mult1_un145_sum_0[1] ));
    NOR2 \d5_RNO[1]  (.A(reset_c), .B(I_12_4), .Y(\d5_RNO[1]_net_1 ));
    DFN1E1 \cur_rand_1[23]  (.D(\d8[2]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[23]));
    AO13 \un2_d5_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I3_CO1  
        (.A(I2_un1_CO1_37), .B(\mult1_un33_sum_0[2] ), .C(
        \mult1_un33_sum_0[4] ), .Y(N89_8));
    XNOR2 \un2_d5_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_11), .B(\mult1_un47_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_34));
    OR2 
        \un2_d6_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I2_un1_CO1_0_tz  
        (.A(\mult1_un166_sum_0[2] ), .B(I1_un3_CO1_2), .Y(
        ADD_5x5_slow_I2_un1_CO1_0_tz_0));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_34), .B(\mult1_un40_sum[2] ), .Y(I3_un3_CO1_6));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_26), .B(\mult1_un75_sum[2] ), .C(
        \mult1_un75_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_35));
    XOR3 \un2_d6_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_S  (
        .A(N83_15), .B(ADD_5x5_slow_I2_S_2), .C(ADD_4x4_slow_I1_S_0), 
        .Y(ADD_5x5_slow_I1_S_0));
    XOR2 \un2_d6_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_0), .B(\mult1_un145_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_0));
    DFN1C0 \rd[9]  (.D(\rd[8]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[9]_net_1 ));
    NOR2A 
        \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_un3_CO1  
        (.A(\rd[0]_net_1 ), .B(\rd[1]_net_1 ), .Y(I1_un3_CO1_6));
    OA1A 
        \un2_d3_if_generate_plus.mult1_un145_sum_ADD_4x4_slow_I1_CO1_0  
        (.A(\rd[5]_net_1 ), .B(\mult1_un138_sum[3] ), .C(\rd[4]_net_1 )
        , .Y(ADD_4x4_slow_I1_CO1_0_1));
    XNOR3 \un2_d5_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un26_sum_0[4] ), .B(\mult1_un26_sum_0[2] ), .C(
        I2_un1_CO1_39), .Y(ADD_5x5_slow_I4_Y_1_14));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_11), .B(\mult1_un82_sum[2] ), .C(
        \mult1_un82_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_0));
    NOR2A 
        \un2_d7_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I1_un2_CO1  
        (.A(\mult1_un159_sum[4] ), .B(\rd[2]_net_1 ), .Y(I1_un2_CO1_6));
    XOR3 \un2_d5_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un68_sum_0[4] ), .B(\mult1_un68_sum_1[1] ), .C(
        N85_30), .Y(\mult1_un75_sum_0[2] ));
    XNOR3 \un2_d3_if_generate_plus.mult1_un96_sum_ADD_4x4_slow_I3_Y_2  
        (.A(N74_10), .B(ADD_4x4_slow_I3_Y_0_5), .C(\mult1_un89_sum[3] )
        , .Y(ADD_4x4_slow_I3_Y_2_9));
    XOR2 \un2_d6_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_2), .B(\mult1_un152_sum[3] ), .Y(
        ADD_5x5_slow_I2_S_1));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_29), .B(\mult1_un61_sum[2] ), .Y(I3_un3_CO1_3));
    XNOR3 
        \un2_d5_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_4), .B(ADD_5x5_slow_I4_Y_0_1), .C(
        \mult1_un166_sum_0[4] ), .Y(ADD_5x5_slow_I4_Y_2_3));
    AO1 \un2_d3_if_generate_plus.mult1_un61_sum_ADD_4x4_slow_I1_CO1  (
        .A(\mult1_un54_sum[3] ), .B(\rd[16]_net_1 ), .C(N74_1_6), .Y(
        N74_14));
    XNOR2 \un2_d7_if_generate_plus.mult1_un19_sum_ADD_5x5_slow_I2_S  (
        .A(N85_0), .B(\rd[23]_net_1 ), .Y(\mult1_un19_sum[2] ));
    AO18 \un2_d5_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un26_sum_0[4] ), .B(\rd[20]_net_1 ), .C(
        \rd[21]_net_1 ), .Y(N85_33));
    XNOR2 \un2_d7_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_12), .B(\mult1_un40_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_35));
    XOR2 \un2_d7_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I4_Y  (
        .A(ADD_5x5_slow_I4_Y_2_33), .B(N89_4), .Y(\mult1_un54_sum[4] ));
    AX1D \un2_d5_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_9), .B(ADD_5x5_slow_I3_CO1_0_8), .C(
        ADD_5x5_slow_I4_Y_2_19), .Y(\mult1_un117_sum_0[4] ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_8), .B(\mult1_un145_sum_0[2] ), .Y(
        I3_un3_CO1_28));
    AX1D \un2_d3_if_generate_plus.mult1_un138_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_4), .B(ADD_4x4_slow_I2_un1_CO1_0_2), .C(
        ADD_4x4_slow_I3_Y_2_3), .Y(\mult1_un138_sum[3] ));
    AO13 \un2_d6_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un131_sum_0[3] ), .B(\rd[6]_net_1 ), .C(
        \rd[7]_net_1 ), .Y(N83_2));
    NOR2 
        \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I1_un2_CO1  
        (.A(\mult1_un75_sum[4] ), .B(\rd[14]_net_1 ), .Y(I1_un2_CO1_10)
        );
    AX1D \un2_d3_if_generate_plus.mult1_un82_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_8), .B(ADD_4x4_slow_I2_un1_CO1_0_6), .C(
        ADD_4x4_slow_I3_Y_2_11), .Y(\mult1_un82_sum[3] ));
    XA1 
        \un2_d6_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I1_un5_CO1  
        (.A(N83_15), .B(ADD_5x5_slow_I2_S_2), .C(\rd[1]_net_1 ), .Y(
        I1_un5_CO1_1));
    XNOR2 \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I1_S  
        (.A(ADD_4x4_slow_I1_S_0_5), .B(\mult1_un117_sum_0[4] ), .Y(
        \mult1_un124_sum_0[1] ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_20), .B(\mult1_un103_sum_0[2] ), .Y(
        I3_un3_CO1_20));
    XNOR2 \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_0), .B(\mult1_un75_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_2));
    NOR2A \d2_RNO_0[0]  (.A(\rd[0]_net_1 ), .B(reset_c), .Y(
        \d2_RNO_0[0]_net_1 ));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un145_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(I1_un3_CO1_4), .B(\mult1_un138_sum_1[1] ), .C(
        \mult1_un138_sum[3] ), .Y(ADD_4x4_slow_I2_un1_CO1_0_3));
    NOR3B 
        \un2_d5_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I2_un5_CO1  
        (.A(\rd[8]_net_1 ), .B(\mult1_un110_sum_0[4] ), .C(
        \rd[9]_net_1 ), .Y(I2_un5_CO1));
    XOR3 \un2_d7_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un117_sum[4] ), .B(\mult1_un117_sum_1[1] ), .C(
        N85_24), .Y(\mult1_un124_sum[2] ));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_0), .B(\mult1_un110_sum_0[2] ), .C(
        \mult1_un110_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_8));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un75_sum_ADD_4x4_slow_I1_CO1_1  
        (.A(\rd[14]_net_1 ), .B(\mult1_un68_sum[3] ), .C(
        \rd[15]_net_1 ), .Y(N74_1_5));
    XNOR2 \un2_d6_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I2_S_2  
        (.A(ADD_5x5_slow_I2_S_1_16), .B(\mult1_un40_sum_1[4] ), .Y(
        ADD_5x5_slow_I2_S_2_16));
    OA1 
        \un2_d5_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(I1_un3_CO1_11), .B(\mult1_un33_sum_1[1] ), .C(
        \mult1_un33_sum_0[4] ), .Y(ADD_5x5_slow_I2_un1_CO1_0_12));
    XNOR2 \un2_d5_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_17), .B(\mult1_un33_sum_0[4] ), .Y(
        \mult1_un40_sum_1[1] ));
    DFN1E1 \cur_rand_1[15]  (.D(\d6[0]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[15]));
    XOR2 \un2_d7_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_13), .B(\mult1_un61_sum[4] ), .Y(
        \mult1_un68_sum_0[1] ));
    OR2 
        \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(ADD_5x5_slow_I2_un1_CO1_0_4), .B(I2_un4_CO1_23), .Y(
        I2_un1_CO1_16));
    XOR2 \un2_d3_if_generate_plus.mult1_un131_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_4), .B(\mult1_un124_sum[3] ), .Y(
        \mult1_un131_sum[1] ));
    AO1 \un2_d7_if_generate_plus.mult1_un1_sum_I_15  (.A(
        \DWACT_ADD_CI_0_pog_array_0[0] ), .B(\DWACT_ADD_CI_0_TMP_0[0] )
        , .C(\DWACT_ADD_CI_0_g_array_0_1[0] ), .Y(
        \DWACT_ADD_CI_0_g_array_1_0[0] ));
    OR2 
        \un2_d7_if_generate_plus.mult1_un19_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\rd[23]_net_1 ), .B(N85_0), .Y(I2_un1_CO1));
    XOR3 \un2_d5_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un40_sum_0[4] ), .B(\mult1_un40_sum_1[1] ), .C(
        N85_28), .Y(\mult1_un47_sum_0[2] ));
    OA1 
        \un2_d5_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(N85_12), .B(\mult1_un19_sum_1[1] ), .C(\mult1_un19_sum[4] )
        , .Y(ADD_5x5_slow_I2_un1_CO1_0_14));
    XA1B 
        \un2_d6_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I1_un2_CO1  
        (.A(N83), .B(ADD_5x5_slow_I2_S_2_0), .C(\rd[3]_net_1 ), .Y(
        I1_un2_CO1_12));
    AO1 
        \un2_d3_if_generate_plus.mult1_un103_sum_ADD_4x4_slow_I2_un1_CO1  
        (.A(N74_8), .B(\mult1_un96_sum[1] ), .C(
        ADD_4x4_slow_I2_un1_CO1_0_13), .Y(I2_un1_CO1_45));
    XOR2 \un2_d3_if_generate_plus.mult1_un82_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_11), .B(\mult1_un75_sum[3] ), .Y(
        \mult1_un82_sum_0[1] ));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_18), .B(\mult1_un152_sum_0[2] ), .C(
        \mult1_un152_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_13));
    NOR2A 
        \un2_d3_if_generate_plus.mult1_un103_sum_ADD_4x4_slow_I2_un1_CO1_0  
        (.A(ADD_4x4_slow_I2_un1_CO1_0_tz_1), .B(\mult1_un96_sum[3] ), 
        .Y(ADD_4x4_slow_I2_un1_CO1_0_13));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_11), .B(\mult1_un124_sum[2] ), .Y(I3_un3_CO1_7));
    AX1D \un2_d5_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_23), .B(ADD_5x5_slow_I3_CO1_0_22), .C(
        ADD_5x5_slow_I4_Y_2_36), .Y(\mult1_un47_sum_0[4] ));
    OR2 
        \un2_d5_if_generate_plus.mult1_un131_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(ADD_5x5_slow_I2_un1_CO1_0_3), .B(I2_un4_CO1_22), .Y(
        I2_un1_CO1_14));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_23), .B(\mult1_un82_sum[2] ), .Y(I3_un3_CO1_1));
    XOR2 \un2_d6_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_5), .B(\mult1_un124_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_3));
    XNOR3 \un2_d5_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un61_sum_0[4] ), .B(\mult1_un61_sum_0[2] ), .C(
        I2_un1_CO1_30), .Y(ADD_5x5_slow_I4_Y_1_6));
    OA1C 
        \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I1_CO1_1  
        (.A(\mult1_un117_sum_0[4] ), .B(\rd[7]_net_1 ), .C(
        \rd[8]_net_1 ), .Y(N85_1_1));
    XOR2 \un2_d6_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_2_11), .B(N83_12), .Y(
        \mult1_un89_sum_0[3] ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(N85_42), .B(\mult1_un82_sum_1[1] ), .Y(I2_un4_CO1_25));
    AO1 
        \un2_d7_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I3_CO1_0_tz  
        (.A(\mult1_un68_sum_0[1] ), .B(N85_5), .C(\mult1_un68_sum[2] ), 
        .Y(ADD_5x5_slow_I3_CO1_0_tz_1));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I1_un5_CO1  
        (.A(\mult1_un82_sum_0[4] ), .B(\rd[12]_net_1 ), .Y(I1_un5_CO1));
    OR2A \un2_d7_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I1_CO1  
        (.A(\rd[22]_net_1 ), .B(\rd[21]_net_1 ), .Y(N85));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_17), .B(\mult1_un145_sum[2] ), .C(
        \mult1_un145_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_15));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_7), .B(\mult1_un131_sum_0[2] ), .C(
        \mult1_un131_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_28));
    OR2 \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I1_CO1  
        (.A(ADD_5x5_slow_I1_CO1_0_3), .B(I1_un2_CO1_8), .Y(N85_21));
    OA1 
        \un2_d5_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(N85_27), .B(\mult1_un110_sum_0[4] ), .C(
        \mult1_un110_sum_1[1] ), .Y(I2_un1_CO1_1_0));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(\mult1_un145_sum_0[1] ), .B(N85_19), .Y(I2_un4_CO1_17));
    XOR2 \un2_d6_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I2_S_1  
        (.A(ADD_4x4_slow_I1_S_0_4), .B(\mult1_un131_sum_0[3] ), .Y(
        ADD_5x5_slow_I2_S_1_2));
    AO13 \un2_d7_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un54_sum[4] ), .B(\rd[16]_net_1 ), .C(
        \rd[17]_net_1 ), .Y(N85_7));
    XOR3 \un2_d5_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un89_sum_0[4] ), .B(\mult1_un89_sum_1[1] ), .C(
        N85_41), .Y(\mult1_un96_sum_0[2] ));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un124_sum_ADD_4x4_slow_I3_Y_2  
        (.A(ADD_4x4_slow_I3_Y_1_3), .B(\mult1_un117_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_2_5));
    AO18 \un2_d6_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I1_CO1  
        (.A(I2_un4_CO1_0), .B(\rd[20]_net_1 ), .C(\rd[21]_net_1 ), .Y(
        N83_13));
    XOR2 \un2_d3_if_generate_plus.mult1_un54_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_15), .B(\mult1_un47_sum[3] ), .Y(
        \mult1_un54_sum[1] ));
    XOR2 \un2_d3_if_generate_plus.mult1_un166_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0), .B(\mult1_un159_sum[3] ), .Y(
        \mult1_un166_sum_0[1] ));
    OR3 \un2_d6_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I1_CO1  
        (.A(I1_un5_CO1_2), .B(I1_un3_CO1_3), .C(I1_un2_CO1_12), .Y(
        N83_15));
    XOR2 \un2_d7_if_generate_plus.mult1_un1_sum_I_12  (.A(
        \DWACT_ADD_CI_0_partial_sum_0[1] ), .B(
        \DWACT_ADD_CI_0_TMP_0[0] ), .Y(I_12_3));
    XNOR3 
        \un2_d5_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_14), .B(ADD_5x5_slow_I4_Y_0_11), .C(
        \mult1_un131_sum_0[4] ), .Y(ADD_5x5_slow_I4_Y_2_13));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un61_sum_ADD_4x4_slow_I1_CO1_1  
        (.A(\rd[16]_net_1 ), .B(\mult1_un54_sum[3] ), .C(
        \rd[17]_net_1 ), .Y(N74_1_6));
    AX1D \un2_d3_if_generate_plus.mult1_un110_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_10), .B(ADD_4x4_slow_I2_un1_CO1_0_8), .C(
        ADD_4x4_slow_I3_Y_2_7), .Y(\mult1_un110_sum[3] ));
    OR2 
        \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I2_un1_CO1_1_tz  
        (.A(N85_2), .B(\mult1_un145_sum[4] ), .Y(I2_un1_CO1_1_tz));
    XOR2 \un2_d7_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_12), .B(\mult1_un68_sum[4] ), .Y(
        \mult1_un75_sum[1] ));
    XOR3 \un2_d7_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un54_sum[4] ), .B(\mult1_un54_sum_0[1] ), .C(N85_7), 
        .Y(\mult1_un61_sum[2] ));
    XNOR2 \un2_d5_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_10), .B(\mult1_un82_sum[4] ), .Y(
        \mult1_un89_sum_1[1] ));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_4), .B(\mult1_un159_sum_0[2] ), .Y(
        I3_un3_CO1_30));
    XNOR2 \un2_d5_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_14), .B(\mult1_un33_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_38));
    XNOR3 
        \un2_d3_if_generate_plus.mult1_un117_sum_ADD_4x4_slow_I3_Y_1  
        (.A(\mult1_un103_sum[3] ), .B(\mult1_un103_sum_0[1] ), .C(
        N74_7), .Y(ADD_4x4_slow_I3_Y_1_4));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_9), .B(\mult1_un103_sum_0[2] ), .C(
        \mult1_un103_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_19));
    XA1B 
        \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I1_un2_CO1  
        (.A(I2_un1_CO1_18), .B(ADD_4x4_slow_I3_Y_2_0), .C(
        \rd[3]_net_1 ), .Y(I1_un2_CO1_14));
    NOR2A 
        \un2_d7_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(ADD_5x5_slow_I3_CO1_0_tz_1), .B(\mult1_un68_sum[4] ), .Y(
        ADD_5x5_slow_I3_CO1_0_3));
    XNOR2 
        \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un145_sum[2] ), .B(\mult1_un145_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_2));
    XNOR3 
        \un2_d7_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I4_Y_2  
        (.A(I2_un1_CO1_11), .B(ADD_5x5_slow_I4_Y_0_8), .C(
        \mult1_un131_sum[4] ), .Y(ADD_5x5_slow_I4_Y_2_10));
    AX1D \un2_d3_if_generate_plus.mult1_un145_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_5), .B(ADD_4x4_slow_I2_un1_CO1_0_3), .C(
        ADD_4x4_slow_I3_Y_2_2), .Y(\mult1_un145_sum[3] ));
    XOR3 \un2_d5_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I2_S  (
        .A(\mult1_un19_sum[4] ), .B(\mult1_un19_sum_1[1] ), .C(N85_12), 
        .Y(\mult1_un26_sum_0[2] ));
    XOR2 \un2_d5_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I4_Y  (
        .A(ADD_5x5_slow_I4_Y_2_30), .B(N89_7), .Y(
        \mult1_un68_sum_0[4] ));
    XOR2 \un2_d3_if_generate_plus.mult1_un68_sum_ADD_4x4_slow_I3_Y  (
        .A(ADD_4x4_slow_I3_Y_2_13), .B(I2_un1_CO1_43), .Y(
        \mult1_un68_sum[3] ));
    AO13 \un2_d7_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I3_CO1  
        (.A(I2_un1_CO1_31), .B(\mult1_un54_sum[2] ), .C(
        \mult1_un54_sum[4] ), .Y(N89_2));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I2_un4_CO1  
        (.A(N85_36), .B(\mult1_un152_sum_1[1] ), .Y(I2_un4_CO1_18));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_3), .B(\mult1_un152_sum[2] ), .Y(I3_un3_CO1_11));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_16), .B(\mult1_un117_sum_0[2] ), .Y(
        I3_un3_CO1_10));
    XNOR2 
        \un2_d7_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un152_sum[2] ), .B(\mult1_un152_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_0));
    AX1D \un2_d5_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I4_Y  (
        .A(I3_un3_CO1_24), .B(ADD_5x5_slow_I3_CO1_0_23), .C(
        ADD_5x5_slow_I4_Y_2_32), .Y(\mult1_un61_sum_0[4] ));
    NOR2B \un2_d5_if_generate_plus.mult1_un1_sum_I_15  (.A(
        \DWACT_ADD_CI_0_TMP[0] ), .B(ADD_5x5_slow_I1_S), .Y(
        \DWACT_ADD_CI_0_g_array_1[0] ));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un166_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[2]_net_1 ), .B(\rd[1]_net_1 ), .Y(ADD_4x4_slow_I1_S_0));
    DFN1C0 \rd[6]  (.D(\rd[5]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[6]_net_1 ));
    OA1 
        \un2_d5_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(I1_un3_CO1_12), .B(\mult1_un26_sum_0[1] ), .C(
        \mult1_un26_sum_0[4] ), .Y(ADD_5x5_slow_I2_un1_CO1_0_13));
    XNOR2 \un2_d3_if_generate_plus.mult1_un47_sum_ADD_4x4_slow_I3_Y_2  
        (.A(ADD_4x4_slow_I3_Y_1_8), .B(\mult1_un40_sum[3] ), .Y(
        ADD_4x4_slow_I3_Y_2_16));
    DFN1C0 \rd[10]  (.D(\rd[9]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[10]_net_1 ));
    OR2 
        \un2_d7_if_generate_plus.mult1_un40_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(ADD_5x5_slow_I2_un1_CO1_0_11), .B(I2_un4_CO1_29), .Y(
        I2_un1_CO1_36));
    NOR2B 
        \un2_d5_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_27), .B(\mult1_un75_sum_0[2] ), .Y(I3_un3_CO1_0)
        );
    NOR3B 
        \un2_d5_if_generate_plus.mult1_un61_sum_ADD_5x5_slow_I2_un5_CO1  
        (.A(\rd[16]_net_1 ), .B(\mult1_un54_sum_0[4] ), .C(
        \rd[17]_net_1 ), .Y(I2_un5_CO1_1));
    DFN1C0 \rd[4]  (.D(\rd[3]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[4]_net_1 ));
    XNOR3 \un2_d7_if_generate_plus.mult1_un54_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un40_sum[4] ), .B(\mult1_un40_sum[2] ), .C(
        I2_un1_CO1_34), .Y(ADD_5x5_slow_I4_Y_1_10));
    MAJ3 
        \un2_d7_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(\mult1_un159_sum[4] ), .B(N85_18), .C(\mult1_un159_sum[1] )
        , .Y(I2_un1_CO1_2));
    XNOR2 
        \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un110_sum_0[2] ), .B(\mult1_un110_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_14));
    OR2 
        \un2_d3_if_generate_plus.mult1_un159_sum_ADD_4x4_slow_I2_un1_CO1_0_tz  
        (.A(\mult1_un152_sum_0[1] ), .B(N74_1_0), .Y(
        ADD_4x4_slow_I2_un1_CO1_0_tz));
    DFN1E1 \cur_rand_1[19]  (.D(\d7[1]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[19]));
    AX1D \un2_d3_if_generate_plus.mult1_un75_sum_ADD_4x4_slow_I3_Y  (
        .A(I2_un4_CO1_2), .B(ADD_4x4_slow_I2_un1_CO1_0_0), .C(
        ADD_4x4_slow_I3_Y_2_12), .Y(\mult1_un75_sum[3] ));
    XOR2 \un2_d7_if_generate_plus.mult1_un33_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_18), .B(\mult1_un26_sum[4] ), .Y(
        \mult1_un33_sum_0[1] ));
    OR2 
        \un2_d5_if_generate_plus.mult1_un145_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(ADD_5x5_slow_I2_un1_CO1_0_2), .B(I2_un4_CO1_20), .Y(
        I2_un1_CO1_10));
    OR2 
        \un2_d3_if_generate_plus.mult1_un103_sum_ADD_4x4_slow_I2_un1_CO1_0_tz  
        (.A(\mult1_un96_sum[1] ), .B(I1_un3_CO1_8), .Y(
        ADD_4x4_slow_I2_un1_CO1_0_tz_1));
    VCC VCC_i (.Y(VCC));
    NOR2A \d5_RNO_0[2]  (.A(I_14_5), .B(reset_c), .Y(
        \d5_RNO_0[2]_net_1 ));
    XNOR2 \un2_d3_if_generate_plus.mult1_un33_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[20]_net_1 ), .B(\rd[21]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_18));
    XNOR2 
        \un2_d5_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I4_Y_2  
        (.A(ADD_5x5_slow_I4_Y_1_5), .B(\mult1_un103_sum_0[4] ), .Y(
        ADD_5x5_slow_I4_Y_2_21));
    DFN1P1C1 \d5[2]  (.D(I_14_5), .CLK(ref_signal_c), .PRE(
        \d5_RNO_0[2]_net_1 ), .CLR(\d5_RNO[2]_net_1 ), .Q(
        \d5[2]_net_1 ));
    XNOR3 
        \un2_d7_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un103_sum[4] ), .B(\mult1_un103_sum[2] ), .C(
        I2_un1_CO1_17), .Y(ADD_5x5_slow_I4_Y_1_2));
    AX1D \un2_d5_if_generate_plus.mult1_un26_sum_ADD_5x5_slow_I4_Y_1  
        (.A(I2_un4_CO1), .B(ADD_5x5_slow_I2_un1_CO1_0), .C(
        \rd[23]_net_1 ), .Y(ADD_5x5_slow_I4_Y_1_16));
    XNOR3 \un2_d7_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I4_Y_1  
        (.A(\mult1_un54_sum[4] ), .B(\mult1_un54_sum[2] ), .C(
        I2_un1_CO1_31), .Y(ADD_5x5_slow_I4_Y_1_7));
    XOR2 \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_1), .B(\mult1_un152_sum[4] ), .Y(
        \mult1_un159_sum[1] ));
    DFN1C0 \rd[0]  (.D(\rd_RNO[0]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[0]_net_1 ));
    AO18 \un2_d5_if_generate_plus.mult1_un68_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un61_sum_0[4] ), .B(\rd[15]_net_1 ), .C(
        \rd[16]_net_1 ), .Y(N85_32));
    OA1B 
        \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un4_CO1_23), .B(\mult1_un117_sum_0[2] ), .C(
        \mult1_un117_sum_0[4] ), .Y(ADD_5x5_slow_I3_CO1_0_9));
    AO13 \un2_d7_if_generate_plus.mult1_un138_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un131_sum[4] ), .B(\rd[5]_net_1 ), .C(\rd[6]_net_1 )
        , .Y(N85_15));
    OR2 
        \un2_d5_if_generate_plus.mult1_un124_sum_ADD_5x5_slow_I2_un1_CO1_0_tz  
        (.A(\mult1_un117_sum_0[1] ), .B(N85_1_1), .Y(
        ADD_5x5_slow_I2_un1_CO1_0_tz));
    XOR2 \un2_d7_if_generate_plus.mult1_un82_sum_ADD_5x5_slow_I2_S  (
        .A(ADD_5x5_slow_I2_S_0_9), .B(N85_3), .Y(\mult1_un82_sum[2] ));
    OR2 
        \un2_d7_if_generate_plus.mult1_un173_sum_ADD_5x5_slow_I2_un1_CO1_1_tz  
        (.A(ADD_5x5_slow_I1_CO1_0_0), .B(\mult1_un166_sum[4] ), .Y(
        I2_un1_CO1_1_tz_1));
    XNOR2 \un2_d5_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un75_sum_0[2] ), .B(\mult1_un75_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_20));
    AO18 \un2_d5_if_generate_plus.mult1_un96_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un89_sum_0[4] ), .B(\rd[11]_net_1 ), .C(
        \rd[12]_net_1 ), .Y(N85_41));
    XOR2 \un2_d7_if_generate_plus.mult1_un89_sum_ADD_5x5_slow_I2_S_0  
        (.A(\mult1_un82_sum[1] ), .B(\mult1_un82_sum_0[4] ), .Y(
        ADD_5x5_slow_I2_S_0_8));
    XNOR3 \un2_d3_if_generate_plus.mult1_un33_sum_ADD_4x4_slow_I3_Y_1  
        (.A(\mult1_un19_sum[3] ), .B(\mult1_un19_sum_0[1] ), .C(N74_19)
        , .Y(ADD_4x4_slow_I3_Y_1_10));
    NOR2A 
        \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I1_un2_CO1  
        (.A(\mult1_un152_sum[4] ), .B(\rd[3]_net_1 ), .Y(I1_un2_CO1_8));
    AO13 \un2_d6_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un110_sum_0[3] ), .B(\rd[9]_net_1 ), .C(
        \rd[10]_net_1 ), .Y(N83_7));
    OR2 \un2_d7_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I1_CO1  
        (.A(ADD_5x5_slow_I1_CO1_0_1), .B(I1_un2_CO1_6), .Y(N85_18));
    XA1 
        \un2_d6_if_generate_plus.mult1_un166_sum_ADD_5x5_slow_I1_un5_CO1  
        (.A(N83), .B(ADD_5x5_slow_I2_S_2_0), .C(\rd[2]_net_1 ), .Y(
        I1_un5_CO1_2));
    XOR2 \un2_d3_if_generate_plus.mult1_un138_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_3), .B(\mult1_un131_sum[3] ), .Y(
        \mult1_un138_sum_1[1] ));
    OA1B 
        \un2_d7_if_generate_plus.mult1_un159_sum_ADD_5x5_slow_I3_CO1_0  
        (.A(I2_un1_CO1_1_4), .B(\mult1_un152_sum[2] ), .C(
        \mult1_un152_sum[4] ), .Y(ADD_5x5_slow_I3_CO1_0_10));
    NOR2A \d7_RNO_0[0]  (.A(\DWACT_ADD_CI_0_partial_sum[0] ), .B(
        reset_c), .Y(\d7_RNO_0[0]_net_1 ));
    XNOR2 
        \un2_d7_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I4_Y_0  
        (.A(\mult1_un138_sum[2] ), .B(\mult1_un138_sum[4] ), .Y(
        ADD_5x5_slow_I4_Y_0_4));
    OA1 
        \un2_d5_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I2_un1_CO1_0  
        (.A(N85_28), .B(\mult1_un40_sum_1[1] ), .C(
        \mult1_un40_sum_0[4] ), .Y(ADD_5x5_slow_I2_un1_CO1_0_10));
    XNOR2 \un2_d3_if_generate_plus.mult1_un75_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[14]_net_1 ), .B(\rd[15]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_12));
    XNOR2 
        \un2_d3_if_generate_plus.mult1_un138_sum_ADD_4x4_slow_I1_S_0  
        (.A(\rd[5]_net_1 ), .B(\rd[6]_net_1 ), .Y(
        ADD_4x4_slow_I1_S_0_3));
    OA1B 
        \un2_d3_if_generate_plus.mult1_un138_sum_ADD_4x4_slow_I1_CO1_1  
        (.A(\mult1_un131_sum[3] ), .B(\rd[5]_net_1 ), .C(\rd[6]_net_1 )
        , .Y(N74_1_1));
    DFN1E1 \cur_rand_1[12]  (.D(\d5[0]_net_1 ), .CLK(ref_signal_c), .E(
        reset_c), .Q(randgen_0_cur_rand[12]));
    XNOR3 
        \un2_d3_if_generate_plus.mult1_un152_sum_ADD_4x4_slow_I3_Y_2  
        (.A(N74_2), .B(ADD_4x4_slow_I3_Y_0_2), .C(\mult1_un145_sum[3] )
        , .Y(ADD_4x4_slow_I3_Y_2_0));
    AO18 \un2_d5_if_generate_plus.mult1_un117_sum_ADD_5x5_slow_I1_CO1  
        (.A(\mult1_un110_sum_0[4] ), .B(\rd[8]_net_1 ), .C(
        \rd[9]_net_1 ), .Y(N85_27));
    NOR2B 
        \un2_d7_if_generate_plus.mult1_un75_sum_ADD_5x5_slow_I3_un3_CO1  
        (.A(I2_un1_CO1_28), .B(\mult1_un68_sum[2] ), .Y(I3_un3_CO1_4));
    XNOR2 \un2_d5_if_generate_plus.mult1_un19_sum_ADD_5x5_slow_I1_S  (
        .A(\rd[22]_net_1 ), .B(\rd[23]_net_1 ), .Y(
        \mult1_un19_sum_1[1] ));
    OR2 \un2_d5_if_generate_plus.mult1_un152_sum_ADD_5x5_slow_I1_CO1  
        (.A(I1_un2_CO1), .B(ADD_5x5_slow_I1_CO1_0), .Y(N85_2));
    XOR2 \un2_d3_if_generate_plus.mult1_un89_sum_ADD_4x4_slow_I1_S  (
        .A(ADD_4x4_slow_I1_S_0_10), .B(\mult1_un82_sum[3] ), .Y(
        \mult1_un89_sum[1] ));
    AO1 
        \un2_d7_if_generate_plus.mult1_un47_sum_ADD_5x5_slow_I2_un1_CO1  
        (.A(N85_11), .B(\mult1_un40_sum[4] ), .C(I2_un1_CO1_1_14), .Y(
        I2_un1_CO1_34));
    OA1 
        \un2_d5_if_generate_plus.mult1_un110_sum_ADD_5x5_slow_I2_un1_CO1_1  
        (.A(N85_40), .B(\mult1_un103_sum_0[4] ), .C(
        \mult1_un103_sum_1[1] ), .Y(I2_un1_CO1_1_9));
    DFN1C0 \rd[7]  (.D(\rd[6]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\rd[7]_net_1 ));
    
endmodule


module two_mhz_clock(
       reset_c,
       GLA,
       clock_out_c
    );
input  reset_c;
input  GLA;
output clock_out_c;

    wire N_11, \counter[1]_net_1 , \counter[0]_net_1 , N_9, 
        \counter[3]_net_1 , \DWACT_FINC_E[0] , N_4, \counter[8]_net_1 , 
        \DWACT_FINC_E[4] , counter14_9, counter14_1, counter14_0, 
        counter14_7, counter14_8, \counter[4]_net_1 , counter14_5, 
        \counter[5]_net_1 , counter14_3, \counter[2]_net_1 , 
        \counter[6]_net_1 , \counter[9]_net_1 , \counter[7]_net_1 , 
        \counter[11]_net_1 , \counter[10]_net_1 , clock_out_RNO_0, 
        \counter_3[5] , I_14_6, \counter_3[4] , I_12_5, \counter_3[1] , 
        I_5_2, I_4_1, I_7_2, I_9_2, I_17_0, I_20_0, I_23_0, I_26_0, 
        I_28, I_32, N_2, \DWACT_FINC_E[6] , \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[5] , N_3, \DWACT_FINC_E[3] , N_5, N_6, N_7, 
        \DWACT_FINC_E[1] , N_8, N_10, GND, VCC;
    
    XOR2 un5_counter_I_5 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .Y(I_5_2));
    XOR2 un5_counter_I_20 (.A(N_6), .B(\counter[7]_net_1 ), .Y(I_20_0));
    NOR2B un5_counter_I_11 (.A(\counter[3]_net_1 ), .B(
        \DWACT_FINC_E[0] ), .Y(N_9));
    XOR2 un5_counter_I_28 (.A(N_3), .B(\counter[10]_net_1 ), .Y(I_28));
    NOR2 \counter_RNIJDL4[11]  (.A(\counter[11]_net_1 ), .B(
        \counter[10]_net_1 ), .Y(counter14_0));
    AND3 un5_counter_I_16 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[1] )
        , .C(\counter[5]_net_1 ), .Y(N_7));
    XOR2 un5_counter_I_17 (.A(N_7), .B(\counter[6]_net_1 ), .Y(I_17_0));
    XOR2 un5_counter_I_32 (.A(N_2), .B(\counter[11]_net_1 ), .Y(I_32));
    AND3 un5_counter_I_29 (.A(\counter[6]_net_1 ), .B(
        \counter[7]_net_1 ), .C(\counter[8]_net_1 ), .Y(
        \DWACT_FINC_E[5] ));
    DFN1C0 \counter[2]  (.D(I_7_2), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[2]_net_1 ));
    DFN1C0 \counter[7]  (.D(I_20_0), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[7]_net_1 ));
    XOR2 un5_counter_I_7 (.A(N_11), .B(\counter[2]_net_1 ), .Y(I_7_2));
    XOR2 un5_counter_I_23 (.A(N_5), .B(\counter[8]_net_1 ), .Y(I_23_0));
    DFN1C0 \counter[6]  (.D(I_17_0), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[6]_net_1 ));
    AOI1B \counter_RNO[4]  (.A(counter14_9), .B(counter14_8), .C(
        I_12_5), .Y(\counter_3[4] ));
    VCC VCC_i (.Y(VCC));
    DFN1C0 \counter[8]  (.D(I_23_0), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[8]_net_1 ));
    AND3 un5_counter_I_22 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\DWACT_FINC_E[3] ), .Y(N_5));
    NOR3C \counter_RNI82AV2[11]  (.A(counter14_1), .B(counter14_0), .C(
        counter14_7), .Y(counter14_9));
    NOR2 \counter_RNI007U[7]  (.A(\counter[9]_net_1 ), .B(
        \counter[7]_net_1 ), .Y(counter14_1));
    AND3 un5_counter_I_8 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(N_10));
    AND3 un5_counter_I_31 (.A(\DWACT_FINC_E[6] ), .B(
        \counter[9]_net_1 ), .C(\counter[10]_net_1 ), .Y(N_2));
    AOI1B \counter_RNO[1]  (.A(counter14_9), .B(counter14_8), .C(I_5_2)
        , .Y(\counter_3[1] ));
    NOR2B un5_counter_I_6 (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(N_11));
    INV un5_counter_I_4 (.A(\counter[0]_net_1 ), .Y(I_4_1));
    AND2 un5_counter_I_15 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(\DWACT_FINC_E[1] ));
    XOR2 un5_counter_I_9 (.A(N_10), .B(\counter[3]_net_1 ), .Y(I_9_2));
    DFN1C0 \counter[4]  (.D(\counter_3[4] ), .CLK(GLA), .CLR(reset_c), 
        .Q(\counter[4]_net_1 ));
    AND2 un5_counter_I_21 (.A(\counter[6]_net_1 ), .B(
        \counter[7]_net_1 ), .Y(\DWACT_FINC_E[3] ));
    DFN1C0 \counter[5]  (.D(\counter_3[5] ), .CLK(GLA), .CLR(reset_c), 
        .Q(\counter[5]_net_1 ));
    XOR2 un5_counter_I_14 (.A(N_8), .B(\counter[5]_net_1 ), .Y(I_14_6));
    XOR2 un5_counter_I_26 (.A(N_4), .B(\counter[9]_net_1 ), .Y(I_26_0));
    AND3 un5_counter_I_27 (.A(\DWACT_FINC_E[4] ), .B(
        \counter[8]_net_1 ), .C(\counter[9]_net_1 ), .Y(N_3));
    AX1C clock_out_RNO (.A(counter14_8), .B(counter14_9), .C(
        clock_out_c), .Y(clock_out_RNO_0));
    AND3 un5_counter_I_10 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(
        \DWACT_FINC_E[0] ));
    GND GND_i (.Y(GND));
    AOI1B \counter_RNO[5]  (.A(counter14_9), .B(counter14_8), .C(
        I_14_6), .Y(\counter_3[5] ));
    AND3 un5_counter_I_18 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .C(\counter[5]_net_1 ), .Y(
        \DWACT_FINC_E[2] ));
    NOR2A \counter_RNIJI6U[0]  (.A(\counter[0]_net_1 ), .B(
        \counter[3]_net_1 ), .Y(counter14_5));
    DFN1C0 \counter[1]  (.D(\counter_3[1] ), .CLK(GLA), .CLR(reset_c), 
        .Q(\counter[1]_net_1 ));
    DFN1C0 \counter[3]  (.D(I_9_2), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[3]_net_1 ));
    AND3 un5_counter_I_19 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\counter[6]_net_1 ), .Y(N_6));
    NOR2 \counter_RNIUT6U[6]  (.A(\counter[8]_net_1 ), .B(
        \counter[6]_net_1 ), .Y(counter14_3));
    NOR3B \counter_RNILKDS1[2]  (.A(\counter[5]_net_1 ), .B(
        counter14_3), .C(\counter[2]_net_1 ), .Y(counter14_7));
    AND3 un5_counter_I_13 (.A(\DWACT_FINC_E[0] ), .B(
        \counter[3]_net_1 ), .C(\counter[4]_net_1 ), .Y(N_8));
    DFN1C0 \counter[11]  (.D(I_32), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[11]_net_1 ));
    XOR2 un5_counter_I_12 (.A(N_9), .B(\counter[4]_net_1 ), .Y(I_12_5));
    AND3 un5_counter_I_30 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\DWACT_FINC_E[5] ), .Y(\DWACT_FINC_E[6] ));
    NOR3B \counter_RNI87DS1[1]  (.A(\counter[4]_net_1 ), .B(
        counter14_5), .C(\counter[1]_net_1 ), .Y(counter14_8));
    NOR2B un5_counter_I_25 (.A(\counter[8]_net_1 ), .B(
        \DWACT_FINC_E[4] ), .Y(N_4));
    DFN1C0 clock_out (.D(clock_out_RNO_0), .CLK(GLA), .CLR(reset_c), 
        .Q(clock_out_c));
    AND3 un5_counter_I_24 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\DWACT_FINC_E[3] ), .Y(\DWACT_FINC_E[4] ));
    DFN1C0 \counter[0]  (.D(I_4_1), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[0]_net_1 ));
    DFN1C0 \counter[10]  (.D(I_28), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[10]_net_1 ));
    DFN1C0 \counter[9]  (.D(I_26_0), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[9]_net_1 ));
    
endmodule


module whitening(
       whitening_0_output_whitening,
       reset_c,
       ref_signal_c,
       data_source_0_output_data,
       output_signal_c
    );
output whitening_0_output_whitening;
input  reset_c;
input  ref_signal_c;
input  data_source_0_output_data;
input  output_signal_c;

    wire N_15, \output_counter[1]_net_1 , \output_counter[0]_net_1 , 
        N_13, \output_counter[3]_net_1 , \DWACT_FINC_E[0] , N_8, 
        \output_counter[8]_net_1 , \DWACT_FINC_E[4] , N_5, 
        \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , counter_n1_i_1, 
        \counter[0]_net_1 , \counter_i_0[1] , counter_n1_i_a3_0_0, 
        \counter[4]_net_1 , \counter[5]_net_1 , state_1_sqmuxa_i_a3_1, 
        output_counter17_13, output_counter17_5, output_counter17_4, 
        output_counter17_11, output_counter17_12, output_counter17_1, 
        output_counter17_0, output_counter17_9, output_counter17_7, 
        \output_counter[12]_net_1 , output_counter17_3, 
        \output_counter[7]_net_1 , \output_counter[2]_net_1 , 
        \output_counter[6]_net_1 , \output_counter[9]_net_1 , 
        \output_counter[4]_net_1 , \output_counter[10]_net_1 , 
        \output_counter[13]_net_1 , \output_counter[5]_net_1 , 
        \output_counter[14]_net_1 , \output_counter[15]_net_1 , 
        \output_counter[11]_net_1 , counter_n5_i_a2_0_9, 
        counter_n5_i_a2_0_6, \counter[14]_net_1 , \counter[9]_net_1 , 
        counter_n5_i_a2_0_8, \counter_i_0[7] , counter_n5_i_a2_0_4, 
        \counter[12]_net_1 , counter_n5_i_a2_0_7, \counter_i_0[2] , 
        counter_n5_i_a2_0_2, \counter[15]_net_1 , \counter_i_0[3] , 
        \counter_i_0[6] , \counter[13]_net_1 , \counter[11]_net_1 , 
        \counter[10]_net_1 , \counter_i_0[8] , output_counter21_13, 
        output_counter21_5, output_counter21_4, output_counter21_11, 
        output_counter21_12, output_counter21_1, output_counter21_9, 
        output_counter21_7, output_whitening_4_i_x2_0, 
        \state[6]_net_1 , N_177, N_11, N_44, N_111, N_13_0, N_42, 
        N_15_0, N_41, N_17, N_114, N_66_i, N_19, N_115, N_65_i, N_21, 
        N_38, N_23, N_37, N_25, output_whitening_1_sqmuxa, 
        \output_counter_5[1] , I_5_3, \output_counter_5[4] , I_12_6, 
        \output_counter_5[5] , I_14_7, \state_22[1] , \state[0]_net_1 , 
        \state_22[2] , \state[1]_net_1 , \state_22[3] , 
        \state[2]_net_1 , \state_22[5] , \state[4]_net_1 , 
        \state_22[6] , \state[5]_net_1 , counter_n0, counter_n15, N_51, 
        counter_n14, N_49, counter_n13, N_48, counter_n12, N_47, 
        counter_n11, N_46, counter_n10, N_45, counter_n9, N_28, 
        \state[3]_net_1 , N_30, N_32, N_34, N_40, I_4_2, I_7_3, I_9_3, 
        I_17_1, I_20_1, I_23_1, I_26_1, I_28_0, I_32_0, I_35_1, I_37_1, 
        I_40_1, I_43, N_2, \DWACT_FINC_E[9] , N_3, \DWACT_FINC_E[8] , 
        N_4, N_6, \DWACT_FINC_E[2] , \DWACT_FINC_E[5] , N_7, 
        \DWACT_FINC_E[3] , N_9, N_10, N_11_0, \DWACT_FINC_E[1] , N_12, 
        N_14, GND, VCC;
    
    DFN1E1C0 \state[0]  (.D(N_30), .CLK(ref_signal_c), .CLR(reset_c), 
        .E(N_34), .Q(\state[0]_net_1 ));
    INV un2_output_counter_1_I_4 (.A(\output_counter[0]_net_1 ), .Y(
        I_4_2));
    NOR2B un2_output_counter_1_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_5));
    DFN0E1C0 \output_counter[14]  (.D(I_40_1), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(output_signal_c), .Q(
        \output_counter[14]_net_1 ));
    DFN0E1C0 \output_counter[13]  (.D(I_37_1), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(output_signal_c), .Q(
        \output_counter[13]_net_1 ));
    NOR2 output_whitening_RNO_7 (.A(\output_counter[14]_net_1 ), .B(
        \output_counter[2]_net_1 ), .Y(output_counter21_1));
    XA1A \counter_RNO[11]  (.A(\counter[11]_net_1 ), .B(N_46), .C(
        output_signal_c), .Y(counter_n11));
    XOR2 un2_output_counter_1_I_37 (.A(N_4), .B(
        \output_counter[13]_net_1 ), .Y(I_37_1));
    DFN0E1C0 \output_counter[5]  (.D(\output_counter_5[5] ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(output_signal_c), .Q(
        \output_counter[5]_net_1 ));
    DFN1C0 \counter[11]  (.D(counter_n11), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[11]_net_1 ));
    NOR3C \output_counter_RNI07MI1[14]  (.A(output_counter17_1), .B(
        output_counter17_0), .C(output_counter17_9), .Y(
        output_counter17_12));
    DFN1E1C0 \state[6]  (.D(\state_22[6] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_34), .Q(\state[6]_net_1 ));
    DFN0E1C0 \output_counter[3]  (.D(I_9_3), .CLK(ref_signal_c), .CLR(
        reset_c), .E(output_signal_c), .Q(\output_counter[3]_net_1 ));
    XOR2 un2_output_counter_1_I_28 (.A(N_7), .B(
        \output_counter[10]_net_1 ), .Y(I_28_0));
    NOR3A \counter_RNIL7DG1[9]  (.A(counter_n5_i_a2_0_6), .B(
        \counter[14]_net_1 ), .C(\counter[9]_net_1 ), .Y(
        counter_n5_i_a2_0_9));
    XA1A \counter_RNO[15]  (.A(\counter[15]_net_1 ), .B(N_51), .C(
        output_signal_c), .Y(counter_n15));
    NOR3A \output_counter_RNIM5IV[2]  (.A(output_counter17_3), .B(
        \output_counter[7]_net_1 ), .C(\output_counter[2]_net_1 ), .Y(
        output_counter17_9));
    AND3 un2_output_counter_1_I_29 (.A(\output_counter[6]_net_1 ), .B(
        \output_counter[7]_net_1 ), .C(\output_counter[8]_net_1 ), .Y(
        \DWACT_FINC_E[5] ));
    NOR3B \counter_RNIJCNS[6]  (.A(\counter_i_0[3] ), .B(
        \counter_i_0[6] ), .C(\counter[13]_net_1 ), .Y(
        counter_n5_i_a2_0_6));
    NOR2 \output_counter_RNIJJ7S[6]  (.A(\output_counter[6]_net_1 ), 
        .B(\output_counter[9]_net_1 ), .Y(output_counter17_5));
    XAI1 \counter_RNO[7]  (.A(N_42), .B(\counter_i_0[7] ), .C(
        output_signal_c), .Y(N_13_0));
    XOR2 un2_output_counter_1_I_43 (.A(N_2), .B(
        \output_counter[15]_net_1 ), .Y(I_43));
    DFN1P0 \counter[6]  (.D(N_15_0), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\counter_i_0[6] ));
    DFN0E1C0 \output_counter[4]  (.D(\output_counter_5[4] ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(output_signal_c), .Q(
        \output_counter[4]_net_1 ));
    XAI1A \counter_RNO_1[1]  (.A(\counter[0]_net_1 ), .B(
        \counter_i_0[1] ), .C(output_signal_c), .Y(counter_n1_i_1));
    DFN1P0 \counter[3]  (.D(N_21), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\counter_i_0[3] ));
    DFN1P0 \counter[2]  (.D(N_23), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\counter_i_0[2] ));
    OR3B \counter_RNO[8]  (.A(output_signal_c), .B(N_44), .C(N_111), 
        .Y(N_11));
    XA1A \counter_RNO[13]  (.A(\counter[13]_net_1 ), .B(N_48), .C(
        output_signal_c), .Y(counter_n13));
    AND3 un2_output_counter_1_I_8 (.A(\output_counter[0]_net_1 ), .B(
        \output_counter[1]_net_1 ), .C(\output_counter[2]_net_1 ), .Y(
        N_14));
    NOR3C \counter_RNO_0[4]  (.A(\counter[0]_net_1 ), .B(
        \counter[5]_net_1 ), .C(N_177), .Y(N_115));
    DFN1E1C0 \state[4]  (.D(N_28), .CLK(ref_signal_c), .CLR(reset_c), 
        .E(N_34), .Q(\state[4]_net_1 ));
    NOR2B un2_output_counter_1_I_11 (.A(\output_counter[3]_net_1 ), .B(
        \DWACT_FINC_E[0] ), .Y(N_13));
    NOR2B un2_output_counter_1_I_6 (.A(\output_counter[1]_net_1 ), .B(
        \output_counter[0]_net_1 ), .Y(N_15));
    XA1A \counter_RNO[12]  (.A(\counter[12]_net_1 ), .B(N_47), .C(
        output_signal_c), .Y(counter_n12));
    AO1 \counter_RNO[1]  (.A(counter_n1_i_a3_0_0), .B(N_177), .C(
        counter_n1_i_1), .Y(N_25));
    NOR3C \counter_RNI3P3V3[9]  (.A(counter_n5_i_a2_0_8), .B(
        counter_n5_i_a2_0_7), .C(counter_n5_i_a2_0_9), .Y(N_177));
    NOR2B \counter_RNO_0[1]  (.A(\counter[4]_net_1 ), .B(
        \counter[5]_net_1 ), .Y(counter_n1_i_a3_0_0));
    NOR2 output_whitening_RNO_5 (.A(\output_counter[1]_net_1 ), .B(
        \output_counter[4]_net_1 ), .Y(output_counter21_4));
    DFN1C0 \counter[4]  (.D(N_19), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[4]_net_1 ));
    DFN1E1C0 \state[5]  (.D(\state_22[5] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_34), .Q(\state[5]_net_1 ));
    DFN1C0 \counter[10]  (.D(counter_n10), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[10]_net_1 ));
    OR2 \counter_RNIPQ4R[2]  (.A(\counter_i_0[2] ), .B(N_37), .Y(N_38));
    GND GND_i (.Y(GND));
    DFN1C0 \counter[13]  (.D(counter_n13), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[13]_net_1 ));
    DFN0E1C0 \output_counter[9]  (.D(I_26_1), .CLK(ref_signal_c), .CLR(
        reset_c), .E(output_signal_c), .Q(\output_counter[9]_net_1 ));
    AND3 un2_output_counter_1_I_33 (.A(\output_counter[9]_net_1 ), .B(
        \output_counter[10]_net_1 ), .C(\output_counter[11]_net_1 ), 
        .Y(\DWACT_FINC_E[7] ));
    DFN1C0 \counter[12]  (.D(counter_n12), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[12]_net_1 ));
    AND3 un2_output_counter_1_I_16 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[1] ), .C(\output_counter[5]_net_1 ), .Y(N_11_0));
    OR2A \counter_RNI8VOF3[11]  (.A(\counter[11]_net_1 ), .B(N_46), .Y(
        N_47));
    NOR2A \output_counter_RNI997S[1]  (.A(\output_counter[4]_net_1 ), 
        .B(\output_counter[1]_net_1 ), .Y(output_counter17_4));
    AND3 un2_output_counter_1_I_42 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[9] ), .Y(N_2));
    NOR3C output_whitening_RNO_2 (.A(output_counter21_1), .B(
        output_counter17_0), .C(output_counter21_9), .Y(
        output_counter21_12));
    AND3 un2_output_counter_1_I_10 (.A(\output_counter[0]_net_1 ), .B(
        \output_counter[1]_net_1 ), .C(\output_counter[2]_net_1 ), .Y(
        \DWACT_FINC_E[0] ));
    NOR3 \counter_RNIV05R[4]  (.A(\counter[5]_net_1 ), .B(
        \counter[4]_net_1 ), .C(\counter[0]_net_1 ), .Y(
        state_1_sqmuxa_i_a3_1));
    XA1 output_whitening_RNO (.A(\state[3]_net_1 ), .B(
        output_whitening_4_i_x2_0), .C(output_signal_c), .Y(N_32));
    NOR3A output_whitening_RNO_8 (.A(output_counter17_3), .B(
        \output_counter[7]_net_1 ), .C(\output_counter[5]_net_1 ), .Y(
        output_counter21_9));
    NOR2B \state_RNO[1]  (.A(\state[0]_net_1 ), .B(output_signal_c), 
        .Y(\state_22[1] ));
    DFN1C0 \counter[15]  (.D(counter_n15), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[15]_net_1 ));
    XOR2 un2_output_counter_1_I_14 (.A(N_12), .B(
        \output_counter[5]_net_1 ), .Y(I_14_7));
    AO1B \counter_RNI4KP75[4]  (.A(state_1_sqmuxa_i_a3_1), .B(N_177), 
        .C(output_signal_c), .Y(N_34));
    OA1 \counter_RNO_0[8]  (.A(N_42), .B(\counter_i_0[7] ), .C(
        \counter_i_0[8] ), .Y(N_111));
    NOR2A \output_counter_RNI777S[0]  (.A(\output_counter[0]_net_1 ), 
        .B(\output_counter[3]_net_1 ), .Y(output_counter17_7));
    VCC VCC_i (.Y(VCC));
    XA1A \counter_RNO[14]  (.A(\counter[14]_net_1 ), .B(N_49), .C(
        output_signal_c), .Y(counter_n14));
    DFN1P0 \counter[1]  (.D(N_25), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\counter_i_0[1] ));
    XOR2 un2_output_counter_1_I_17 (.A(N_11_0), .B(
        \output_counter[6]_net_1 ), .Y(I_17_1));
    NOR3A \counter_RNO[5]  (.A(output_signal_c), .B(N_114), .C(N_66_i), 
        .Y(N_17));
    AND2 un2_output_counter_1_I_21 (.A(\output_counter[6]_net_1 ), .B(
        \output_counter[7]_net_1 ), .Y(\DWACT_FINC_E[3] ));
    NOR2B \state_RNO[4]  (.A(\state[3]_net_1 ), .B(output_signal_c), 
        .Y(N_28));
    XAI1 \counter_RNO[3]  (.A(N_38), .B(\counter_i_0[3] ), .C(
        output_signal_c), .Y(N_21));
    XOR2 un2_output_counter_1_I_32 (.A(N_6), .B(
        \output_counter[11]_net_1 ), .Y(I_32_0));
    OR2A \counter_RNIJQ054[13]  (.A(\counter[13]_net_1 ), .B(N_48), .Y(
        N_49));
    XOR2 un2_output_counter_1_I_35 (.A(N_5), .B(
        \output_counter[12]_net_1 ), .Y(I_35_1));
    NOR2B \state_RNO[2]  (.A(\state[1]_net_1 ), .B(output_signal_c), 
        .Y(\state_22[2] ));
    DFN1C0 \counter[5]  (.D(N_17), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[5]_net_1 ));
    DFN0E1C0 \output_counter[12]  (.D(I_35_1), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(output_signal_c), .Q(
        \output_counter[12]_net_1 ));
    XA1A \counter_RNO[10]  (.A(\counter[10]_net_1 ), .B(N_45), .C(
        output_signal_c), .Y(counter_n10));
    NOR2B \counter_RNIDE3I[1]  (.A(\counter_i_0[1] ), .B(
        \counter_i_0[8] ), .Y(counter_n5_i_a2_0_2));
    XOR2 un2_output_counter_1_I_26 (.A(N_8), .B(
        \output_counter[9]_net_1 ), .Y(I_26_1));
    NOR2B \state_RNO[6]  (.A(\state[5]_net_1 ), .B(output_signal_c), 
        .Y(\state_22[6] ));
    DFN0E1C0 \output_counter[1]  (.D(\output_counter_5[1] ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(output_signal_c), .Q(
        \output_counter[1]_net_1 ));
    XOR2 output_whitening_RNO_3 (.A(\state[6]_net_1 ), .B(
        data_source_0_output_data), .Y(output_whitening_4_i_x2_0));
    NOR3C \counter_RNO_0[5]  (.A(\counter[0]_net_1 ), .B(
        \counter[4]_net_1 ), .C(N_177), .Y(N_114));
    XOR2 un2_output_counter_1_I_20 (.A(N_10), .B(
        \output_counter[7]_net_1 ), .Y(I_20_1));
    OR2 \counter_RNIJNBV1[6]  (.A(N_41), .B(\counter_i_0[6] ), .Y(N_42)
        );
    NOR3B \counter_RNI93P51[15]  (.A(\counter_i_0[2] ), .B(
        counter_n5_i_a2_0_2), .C(\counter[15]_net_1 ), .Y(
        counter_n5_i_a2_0_7));
    AOI1B \output_counter_RNO[1]  (.A(output_counter17_13), .B(
        output_counter17_12), .C(I_5_3), .Y(\output_counter_5[1] ));
    XAI1 \counter_RNO[6]  (.A(\counter_i_0[6] ), .B(N_41), .C(
        output_signal_c), .Y(N_15_0));
    AND3 un2_output_counter_1_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E[4] ));
    OR2A \counter_RNI18HQ2[9]  (.A(\counter[9]_net_1 ), .B(N_44), .Y(
        N_45));
    NOR3A \output_counter_RNI6E0C1[12]  (.A(output_counter17_7), .B(
        \output_counter[12]_net_1 ), .C(\output_counter[8]_net_1 ), .Y(
        output_counter17_11));
    XOR2 un2_output_counter_1_I_5 (.A(\output_counter[0]_net_1 ), .B(
        \output_counter[1]_net_1 ), .Y(I_5_3));
    AND3 un2_output_counter_1_I_13 (.A(\DWACT_FINC_E[0] ), .B(
        \output_counter[3]_net_1 ), .C(\output_counter[4]_net_1 ), .Y(
        N_12));
    AND2 un2_output_counter_1_I_38 (.A(\output_counter[12]_net_1 ), .B(
        \output_counter[13]_net_1 ), .Y(\DWACT_FINC_E[8] ));
    AND3 un2_output_counter_1_I_27 (.A(\DWACT_FINC_E[4] ), .B(
        \output_counter[8]_net_1 ), .C(\output_counter[9]_net_1 ), .Y(
        N_7));
    DFN1E1C0 \state[3]  (.D(\state_22[3] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_34), .Q(\state[3]_net_1 ));
    AND3 un2_output_counter_1_I_39 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[8] ), .Y(N_3));
    NOR3A output_whitening_RNO_6 (.A(output_counter21_7), .B(
        \output_counter[12]_net_1 ), .C(\output_counter[9]_net_1 ), .Y(
        output_counter21_11));
    DFN1C0 \counter[14]  (.D(counter_n14), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[14]_net_1 ));
    AX1D \counter_RNO_1[4]  (.A(N_38), .B(\counter_i_0[3] ), .C(
        \counter[4]_net_1 ), .Y(N_65_i));
    OR2A \counter_RNI563I[1]  (.A(\counter[0]_net_1 ), .B(
        \counter_i_0[1] ), .Y(N_37));
    NOR3B \counter_RNI5ET81[12]  (.A(\counter_i_0[7] ), .B(
        counter_n5_i_a2_0_4), .C(\counter[12]_net_1 ), .Y(
        counter_n5_i_a2_0_8));
    DFN0E1C0 \output_counter[8]  (.D(I_23_1), .CLK(ref_signal_c), .CLR(
        reset_c), .E(output_signal_c), .Q(\output_counter[8]_net_1 ));
    XOR2 \counter_RNO_1[5]  (.A(N_40), .B(\counter[5]_net_1 ), .Y(
        N_66_i));
    NOR3C \output_counter_RNI2BF43[12]  (.A(output_counter17_5), .B(
        output_counter17_4), .C(output_counter17_11), .Y(
        output_counter17_13));
    DFN0E1C0 \output_counter[0]  (.D(I_4_2), .CLK(ref_signal_c), .CLR(
        reset_c), .E(output_signal_c), .Q(\output_counter[0]_net_1 ));
    NOR3A \counter_RNO[4]  (.A(output_signal_c), .B(N_115), .C(N_65_i), 
        .Y(N_19));
    XOR2 un2_output_counter_1_I_7 (.A(N_15), .B(
        \output_counter[2]_net_1 ), .Y(I_7_3));
    NOR2B \state_RNO[5]  (.A(\state[4]_net_1 ), .B(output_signal_c), 
        .Y(\state_22[5] ));
    XOR2 un2_output_counter_1_I_12 (.A(N_13), .B(
        \output_counter[4]_net_1 ), .Y(I_12_6));
    AND2 un2_output_counter_1_I_15 (.A(\output_counter[3]_net_1 ), .B(
        \output_counter[4]_net_1 ), .Y(\DWACT_FINC_E[1] ));
    NOR2 output_whitening_RNO_4 (.A(\output_counter[6]_net_1 ), .B(
        \output_counter[8]_net_1 ), .Y(output_counter21_5));
    DFN1E1C0 \state[2]  (.D(\state_22[2] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_34), .Q(\state[2]_net_1 ));
    AND3 un2_output_counter_1_I_41 (.A(\output_counter[12]_net_1 ), .B(
        \output_counter[13]_net_1 ), .C(\output_counter[14]_net_1 ), 
        .Y(\DWACT_FINC_E[9] ));
    DFN0E1C0 \output_counter[11]  (.D(I_32_0), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(output_signal_c), .Q(
        \output_counter[11]_net_1 ));
    XOR2 un2_output_counter_1_I_23 (.A(N_9), .B(
        \output_counter[8]_net_1 ), .Y(I_23_1));
    NOR2A \output_counter_RNIU5PF[14]  (.A(\output_counter[5]_net_1 ), 
        .B(\output_counter[14]_net_1 ), .Y(output_counter17_1));
    DFN1E1C0 \state[1]  (.D(\state_22[1] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_34), .Q(\state[1]_net_1 ));
    DFN0E1C0 \output_counter[10]  (.D(I_28_0), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(output_signal_c), .Q(
        \output_counter[10]_net_1 ));
    DFN1P0 \counter[7]  (.D(N_13_0), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\counter_i_0[7] ));
    NOR2 output_whitening_RNO_9 (.A(\output_counter[3]_net_1 ), .B(
        \output_counter[0]_net_1 ), .Y(output_counter21_7));
    OR2A \counter_RNIRU9M1[5]  (.A(\counter[5]_net_1 ), .B(N_40), .Y(
        N_41));
    DFN0E1C0 \output_counter[7]  (.D(I_20_1), .CLK(ref_signal_c), .CLR(
        reset_c), .E(output_signal_c), .Q(\output_counter[7]_net_1 ));
    DFN0E0C0 output_whitening (.D(N_32), .CLK(ref_signal_c), .CLR(
        reset_c), .E(output_whitening_1_sqmuxa), .Q(
        whitening_0_output_whitening));
    OR2A \counter_RNO_0[15]  (.A(\counter[14]_net_1 ), .B(N_49), .Y(
        N_51));
    NOR2A \counter_RNO[0]  (.A(output_signal_c), .B(\counter[0]_net_1 )
        , .Y(counter_n0));
    NOR2 \output_counter_RNI9OA3[10]  (.A(\output_counter[10]_net_1 ), 
        .B(\output_counter[13]_net_1 ), .Y(output_counter17_3));
    NOR2B \state_RNO[3]  (.A(\state[2]_net_1 ), .B(output_signal_c), 
        .Y(\state_22[3] ));
    NOR2B \state_RNO[0]  (.A(data_source_0_output_data), .B(
        output_signal_c), .Y(N_30));
    OR3A \counter_RNI478D1[3]  (.A(\counter[4]_net_1 ), .B(N_38), .C(
        \counter_i_0[3] ), .Y(N_40));
    OR3 \counter_RNI6CFH2[8]  (.A(N_42), .B(\counter_i_0[7] ), .C(
        \counter_i_0[8] ), .Y(N_44));
    DFN0E1C0 \output_counter[15]  (.D(I_43), .CLK(ref_signal_c), .CLR(
        reset_c), .E(output_signal_c), .Q(\output_counter[15]_net_1 ));
    XOR2 un2_output_counter_1_I_40 (.A(N_3), .B(
        \output_counter[14]_net_1 ), .Y(I_40_1));
    NOR2 \output_counter_RNICRA3[15]  (.A(\output_counter[15]_net_1 ), 
        .B(\output_counter[11]_net_1 ), .Y(output_counter17_0));
    NOR2 \counter_RNI7N7L[10]  (.A(\counter[11]_net_1 ), .B(
        \counter[10]_net_1 ), .Y(counter_n5_i_a2_0_4));
    AOI1B \output_counter_RNO[4]  (.A(output_counter17_13), .B(
        output_counter17_12), .C(I_12_6), .Y(\output_counter_5[4] ));
    AOI1B \output_counter_RNO[5]  (.A(output_counter17_13), .B(
        output_counter17_12), .C(I_14_7), .Y(\output_counter_5[5] ));
    AND3 un2_output_counter_1_I_31 (.A(\DWACT_FINC_E[6] ), .B(
        \output_counter[9]_net_1 ), .C(\output_counter[10]_net_1 ), .Y(
        N_6));
    AND3 un2_output_counter_1_I_18 (.A(\output_counter[3]_net_1 ), .B(
        \output_counter[4]_net_1 ), .C(\output_counter[5]_net_1 ), .Y(
        \DWACT_FINC_E[2] ));
    AND3 un2_output_counter_1_I_19 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\output_counter[6]_net_1 ), .Y(N_10));
    AOI1B output_whitening_RNO_0 (.A(output_counter21_13), .B(
        output_counter21_12), .C(output_signal_c), .Y(
        output_whitening_1_sqmuxa));
    XAI1 \counter_RNO[2]  (.A(N_37), .B(\counter_i_0[2] ), .C(
        output_signal_c), .Y(N_23));
    DFN1C0 \counter[9]  (.D(counter_n9), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[9]_net_1 ));
    AND3 un2_output_counter_1_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_9));
    OR2A \counter_RNIDSCQ3[12]  (.A(\counter[12]_net_1 ), .B(N_47), .Y(
        N_48));
    NOR2B un2_output_counter_1_I_25 (.A(\output_counter[8]_net_1 ), .B(
        \DWACT_FINC_E[4] ), .Y(N_8));
    XA1A \counter_RNO[9]  (.A(\counter[9]_net_1 ), .B(N_44), .C(
        output_signal_c), .Y(counter_n9));
    AND3 un2_output_counter_1_I_36 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\output_counter[12]_net_1 ), .Y(N_4));
    DFN1P0 \counter[8]  (.D(N_11), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\counter_i_0[8] ));
    XOR2 un2_output_counter_1_I_9 (.A(N_14), .B(
        \output_counter[3]_net_1 ), .Y(I_9_3));
    OR2A \counter_RNI43553[10]  (.A(\counter[10]_net_1 ), .B(N_45), .Y(
        N_46));
    AND3 un2_output_counter_1_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[6] ));
    DFN1C0 \counter[0]  (.D(counter_n0), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[0]_net_1 ));
    DFN0E1C0 \output_counter[2]  (.D(I_7_3), .CLK(ref_signal_c), .CLR(
        reset_c), .E(output_signal_c), .Q(\output_counter[2]_net_1 ));
    NOR3C output_whitening_RNO_1 (.A(output_counter21_5), .B(
        output_counter21_4), .C(output_counter21_11), .Y(
        output_counter21_13));
    DFN0E1C0 \output_counter[6]  (.D(I_17_1), .CLK(ref_signal_c), .CLR(
        reset_c), .E(output_signal_c), .Q(\output_counter[6]_net_1 ));
    
endmodule


module main_clock(
       reset_c,
       GLA,
       ref_signal_c
    );
input  reset_c;
input  GLA;
output ref_signal_c;

    wire clock_out_i, N_7, \counter[1]_net_1 , \counter[0]_net_1 , N_5, 
        \counter[3]_net_1 , \DWACT_FINC_E[0] , counter14_4, 
        counter14_2, \counter[2]_net_1 , \counter[5]_net_1 , 
        counter14_3, \counter[6]_net_1 , \counter[7]_net_1 , 
        \counter[4]_net_1 , clock_out_RNO_net_1, \counter_3[0] , I_5_1, 
        I_7_1, I_9_1, I_12_2, I_14_2, I_17, I_20, N_2, 
        \DWACT_FINC_E[2] , N_3, \DWACT_FINC_E[1] , N_4, N_6, GND, VCC;
    
    NOR2B un5_counter_1_I_11 (.A(\counter[3]_net_1 ), .B(
        \DWACT_FINC_E[0] ), .Y(N_5));
    DFN1C0 \counter[2]  (.D(I_7_1), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[2]_net_1 ));
    DFN1C0 \counter[7]  (.D(I_20), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[7]_net_1 ));
    AND3 un5_counter_1_I_19 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\counter[6]_net_1 ), .Y(N_2));
    XOR2 un5_counter_1_I_12 (.A(N_5), .B(\counter[4]_net_1 ), .Y(
        I_12_2));
    AOI1 \counter_RNO[0]  (.A(counter14_4), .B(counter14_3), .C(
        \counter[0]_net_1 ), .Y(\counter_3[0] ));
    DFN1C0 \counter[6]  (.D(I_17), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[6]_net_1 ));
    VCC VCC_i (.Y(VCC));
    AND3 un5_counter_1_I_18 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .C(\counter[5]_net_1 ), .Y(
        \DWACT_FINC_E[2] ));
    AND3 un5_counter_1_I_10 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(
        \DWACT_FINC_E[0] ));
    XOR2 un5_counter_1_I_9 (.A(N_6), .B(\counter[3]_net_1 ), .Y(I_9_1));
    AND3 un5_counter_1_I_8 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(N_6));
    NOR2B un5_counter_1_I_6 (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(N_7));
    AND3 un5_counter_1_I_13 (.A(\DWACT_FINC_E[0] ), .B(
        \counter[3]_net_1 ), .C(\counter[4]_net_1 ), .Y(N_4));
    DFN1C0 \counter[4]  (.D(I_12_2), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[4]_net_1 ));
    XOR2 un5_counter_1_I_20 (.A(N_2), .B(\counter[7]_net_1 ), .Y(I_20));
    DFN1C0 \counter[5]  (.D(I_14_2), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[5]_net_1 ));
    XOR2 un5_counter_1_I_14 (.A(N_4), .B(\counter[5]_net_1 ), .Y(
        I_14_2));
    XOR2 un5_counter_1_I_7 (.A(N_7), .B(\counter[2]_net_1 ), .Y(I_7_1));
    XOR2 un5_counter_1_I_17 (.A(N_3), .B(\counter[6]_net_1 ), .Y(I_17));
    AND3 un5_counter_1_I_16 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[1] ), .C(\counter[5]_net_1 ), .Y(N_3));
    AX1C clock_out_RNO (.A(counter14_3), .B(counter14_4), .C(
        clock_out_i), .Y(clock_out_RNO_net_1));
    GND GND_i (.Y(GND));
    DFN1C0 \counter[1]  (.D(I_5_1), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[1]_net_1 ));
    CLKINT clock_out_RNIG44 (.A(clock_out_i), .Y(ref_signal_c));
    DFN1C0 \counter[3]  (.D(I_9_1), .CLK(GLA), .CLR(reset_c), .Q(
        \counter[3]_net_1 ));
    XOR2 un5_counter_1_I_5 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .Y(I_5_1));
    NOR3 \counter_RNIFVEB1[7]  (.A(\counter[6]_net_1 ), .B(
        \counter[7]_net_1 ), .C(\counter[3]_net_1 ), .Y(counter14_3));
    NOR2 \counter_RNIF4VS[1]  (.A(\counter[4]_net_1 ), .B(
        \counter[1]_net_1 ), .Y(counter14_2));
    NOR3A \counter_RNI0BUP1[2]  (.A(counter14_2), .B(
        \counter[2]_net_1 ), .C(\counter[5]_net_1 ), .Y(counter14_4));
    AND2 un5_counter_1_I_15 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(\DWACT_FINC_E[1] ));
    DFN1C0 clock_out (.D(clock_out_RNO_net_1), .CLK(GLA), .CLR(reset_c)
        , .Q(clock_out_i));
    DFN1C0 \counter[0]  (.D(\counter_3[0] ), .CLK(GLA), .CLR(reset_c), 
        .Q(\counter[0]_net_1 ));
    
endmodule


module pll_core(
       clock_c,
       GLA
    );
input  clock_c;
output GLA;

    wire CLKAP, Core_GLB, Core_GLC, LOCK, Core_YB, Core_YC, 
        pll_core_GND, pll_core_VCC;
    
    PLL #( .VCOFREQUENCY(100.000000) )  Core (.CLKA(CLKAP), .EXTFB(
        pll_core_GND), .POWERDOWN(pll_core_VCC), .GLA(GLA), .LOCK(LOCK)
        , .GLB(Core_GLB), .YB(Core_YB), .GLC(Core_GLC), .YC(Core_YC), 
        .OADIV0(pll_core_GND), .OADIV1(pll_core_GND), .OADIV2(
        pll_core_GND), .OADIV3(pll_core_GND), .OADIV4(pll_core_GND), 
        .OAMUX0(pll_core_GND), .OAMUX1(pll_core_GND), .OAMUX2(
        pll_core_VCC), .DLYGLA0(pll_core_GND), .DLYGLA1(pll_core_GND), 
        .DLYGLA2(pll_core_GND), .DLYGLA3(pll_core_GND), .DLYGLA4(
        pll_core_GND), .OBDIV0(pll_core_GND), .OBDIV1(pll_core_GND), 
        .OBDIV2(pll_core_GND), .OBDIV3(pll_core_GND), .OBDIV4(
        pll_core_GND), .OBMUX0(pll_core_GND), .OBMUX1(pll_core_GND), 
        .OBMUX2(pll_core_GND), .DLYYB0(pll_core_GND), .DLYYB1(
        pll_core_GND), .DLYYB2(pll_core_GND), .DLYYB3(pll_core_GND), 
        .DLYYB4(pll_core_GND), .DLYGLB0(pll_core_GND), .DLYGLB1(
        pll_core_GND), .DLYGLB2(pll_core_GND), .DLYGLB3(pll_core_GND), 
        .DLYGLB4(pll_core_GND), .OCDIV0(pll_core_GND), .OCDIV1(
        pll_core_GND), .OCDIV2(pll_core_GND), .OCDIV3(pll_core_GND), 
        .OCDIV4(pll_core_GND), .OCMUX0(pll_core_GND), .OCMUX1(
        pll_core_GND), .OCMUX2(pll_core_GND), .DLYYC0(pll_core_GND), 
        .DLYYC1(pll_core_GND), .DLYYC2(pll_core_GND), .DLYYC3(
        pll_core_GND), .DLYYC4(pll_core_GND), .DLYGLC0(pll_core_GND), 
        .DLYGLC1(pll_core_GND), .DLYGLC2(pll_core_GND), .DLYGLC3(
        pll_core_GND), .DLYGLC4(pll_core_GND), .FINDIV0(pll_core_VCC), 
        .FINDIV1(pll_core_VCC), .FINDIV2(pll_core_GND), .FINDIV3(
        pll_core_GND), .FINDIV4(pll_core_GND), .FINDIV5(pll_core_GND), 
        .FINDIV6(pll_core_GND), .FBDIV0(pll_core_VCC), .FBDIV1(
        pll_core_VCC), .FBDIV2(pll_core_GND), .FBDIV3(pll_core_GND), 
        .FBDIV4(pll_core_VCC), .FBDIV5(pll_core_GND), .FBDIV6(
        pll_core_GND), .FBDLY0(pll_core_GND), .FBDLY1(pll_core_GND), 
        .FBDLY2(pll_core_GND), .FBDLY3(pll_core_GND), .FBDLY4(
        pll_core_GND), .FBSEL0(pll_core_VCC), .FBSEL1(pll_core_GND), 
        .XDLYSEL(pll_core_GND), .VCOSEL0(pll_core_GND), .VCOSEL1(
        pll_core_GND), .VCOSEL2(pll_core_VCC));
    PLLINT pllint1 (.A(clock_c), .Y(CLKAP));
    VCC VCC_i (.Y(pll_core_VCC));
    GND GND_i (.Y(pll_core_GND));
    
endmodule


module mac(
       demodulator_0_cur_flag,
       demodulator_0_cur_scheme,
       randgen_0_cur_rand,
       demodulator_0_ord,
       demodulator_0_ctg,
       mac_0_datacmd,
       mac_0_head,
       mac_0_working,
       mac_0_sending,
       reset_c,
       ref_signal_c
    );
input  [7:0] demodulator_0_cur_flag;
input  [47:0] demodulator_0_cur_scheme;
input  [23:3] randgen_0_cur_rand;
input  [1:0] demodulator_0_ord;
input  [1:0] demodulator_0_ctg;
output mac_0_datacmd;
output mac_0_head;
output mac_0_working;
output mac_0_sending;
input  reset_c;
input  ref_signal_c;

    wire init_2_net_1, N_42, init_1_net_1, init_0_net_1, 
        un1_start_1_sqmuxa_3_0, N_401, start_1_sqmuxa, N_400, 
        \DWACT_ADD_CI_0_g_array_11[0] , \DWACT_ADD_CI_0_g_array_2[0] , 
        \DWACT_ADD_CI_0_pog_array_1_1[0] , 
        \DWACT_ADD_CI_0_g_array_3[0] , \DWACT_ADD_CI_0_pog_array_2[0] , 
        \DWACT_ADD_CI_0_g_array_1[0] , \DWACT_ADD_CI_0_pog_array_1[0] , 
        \DWACT_ADD_CI_0_g_array_11_0[0] , 
        \DWACT_ADD_CI_0_g_array_2_0[0] , 
        \DWACT_ADD_CI_0_pog_array_1_1_0[0] , 
        \DWACT_ADD_CI_0_g_array_3_0[0] , 
        \DWACT_ADD_CI_0_pog_array_2_0[0] , 
        \DWACT_ADD_CI_0_g_array_1_0[0] , 
        \DWACT_ADD_CI_0_pog_array_1_0[0] , 
        \DWACT_ADD_CI_0_g_array_12_3[0] , \tick[8]_net_1 , 
        \DWACT_ADD_CI_0_g_array_12[0] , \tick[2]_net_1 , 
        \DWACT_ADD_CI_0_g_array_12_1[0] , \tick[4]_net_1 , 
        \DWACT_ADD_CI_0_g_array_12_2[0] , \tick[6]_net_1 , 
        \DWACT_ADD_CI_0_TMP[0] , \tick[1]_net_1 , 
        \DWACT_ADD_CI_0_g_array_12_3_0[0] , \counter[8]_net_1 , 
        \DWACT_ADD_CI_0_g_array_12_0[0] , \counter[2]_net_1 , 
        \DWACT_ADD_CI_0_g_array_12_1_0[0] , \counter[4]_net_1 , 
        \DWACT_ADD_CI_0_g_array_12_2_0[0] , \counter[6]_net_1 , 
        \DWACT_ADD_CI_0_TMP_0[0] , \counter[1]_net_1 , N_5, 
        \div_counter[1]_net_1 , \div_counter[0]_net_1 , N_3, 
        \div_counter[3]_net_1 , \DWACT_FINC_E[0] , 
        sending_7_i_i_a3_1_0_net_1, memo26, N_329, N_407, N_884, N_312, 
        N_354, ADD_10x10_slow_I8_S_0, \frame_begin[8]_net_1 , 
        \un1_choice_2[8] , ADD_10x10_slow_I7_S_0, 
        \frame_begin[7]_net_1 , \un1_choice_2[7] , 
        \frame_begin_18_i_0_0[6] , \choice[2]_net_1 , N_284, N_505, 
        cnt_n3_0, \cnt[3]_net_1 , cnt_0_sqmuxa, un1_start_1_sqmuxa_5, 
        \frame_begin_18_i_0_0[5] , \choice[1]_net_1 , cnt_n2_0, 
        \cnt[2]_net_1 , \frame_begin_18_i_0_0[4] , N_514, 
        \tick_14_0_0_o2_2[4] , start_net_1, N_296, un1_tick_2_sqmuxa_2, 
        \tick_14_0_0_o2_1[4] , N_314, N_249, N_461, 
        un1_tick_2_sqmuxa_0, start_0_sqmuxa, un1_tick_2_sqmuxa_10_1, 
        N_506, un1_tick_2_sqmuxa_5, un1_calculating_0_sqmuxa_0_0_0, 
        un1_calculating_0_sqmuxa_0_0_a3_0, N_482, 
        un1_resuming_0_sqmuxa_5_0_0_0, N_385, N_371, rd_0_sqmuxa_1_1, 
        \rd[0]_net_1 , \rd[2]_net_1 , \rd[1]_net_1 , 
        ADD_10x10_slow_I3_S_0, \frame_begin[3]_net_1 , I2_un1_CO1, 
        un1_start_1_sqmuxa_7_0_1_0, N_479, N_481, 
        resuming_0_sqmuxa_2_0_a2_0_a3_2, 
        resuming_0_sqmuxa_2_0_a2_0_a3_1, \cnt[1]_net_1 , 
        \cnt[0]_net_1 , un1_start_1_sqmuxa_4_0, tick_2_sqmuxa, 
        ilde_0_0_0, un1_i44, un1_start_1_sqmuxa_1_0_0_0, 
        un1_start_1_sqmuxa_1_0_0_a3_0, N_443, cnt_0_sqmuxa_0, N_259, 
        \flag[0]_net_1 , rd_0_sqmuxa_0, calculating_net_1, N_277, 
        \un1_choice_2_0_a2_0[3] , un1_resuming_0_sqmuxa_5_0_0_o2_0, 
        un1_resuming_0_sqmuxa_5_0_0_o2_1, counting_net_1, 
        tick_1_sqmuxa_2_i_i_o2_0, un1_tick_2_sqmuxa_5_0_0, blank18, 
        start_2_sqmuxa, N_154, head_13_0_i_0, N_361, N_245, N_384, 
        tick_1_sqmuxa_3_i_i_a3_0, resuming_net_1, tick_2_sqmuxa_1, 
        N_274, \tick_14_0_0_a3_2_2_0[4] , N_252, N_449, 
        awaitbeacon_net_1, N_472, choosing_net_1, sending_7_i_i_0, 
        sending_7_i_i_a3_0_0, N_276, data_size_1_sqmuxa_i_0_0, N_288, 
        N_478, un1_tick_1_sqmuxa_2_i_i_a3_1, div_counter11, 
        sending_7_i_i_a3_2_0, launch_net_1, un1_tick_2_sqmuxa_5_0_a2_3, 
        un1_tick_2_sqmuxa_5_0_a2_1, past_net_1, N_264, 
        un1_tick_0_sqmuxa_1_0_0_0_0, N_477, N_480, N_291, 
        id_1_sqmuxa_1_i_0_0, N_292, sending_7_i_i_o2_0_1, N_465, 
        blank_net_1, N_509, start_2_sqmuxa_0, 
        un1_start_0_sqmuxa_0_0_a3_1, N_476, N_263, 
        un1_resuming_0_sqmuxa_5_0_0_a3_1, init_net_1, 
        awaitbeacon_0_i_a3_0, N_309, awaitscheme_6_0_0_o2_0, 
        awaitscheme_6_0_0_o2_4_0, awaitscheme_6_0_0_o2_4_1, N_281, 
        awaitscheme_6_0_0_a3_0_0, N_500, awaitheartbeat_net_1, 
        un1_resuming_0_sqmuxa_5_0_0_a2_0, memo_0_sqmuxa_1_i_i_a3_0, 
        N_501, id_1_sqmuxa_1_i_0_a2_0, \tick[0]_net_1 , 
        un1_start_0_sqmuxa_0_0_a2_0_0, sending13, div_counter11_2, 
        div_counter11_1, \div_counter[2]_net_1 , div_counter11_0, 
        \div_counter[5]_net_1 , \div_counter[4]_net_1 , 
        un1_resuming_0_sqmuxa_3_0_0_o3_0, \i[3]_net_1 , \i[2]_net_1 , 
        un1_tick_0_sqmuxa_1_0_0_o2_1, blank17_NE_6, blank17_NE_0, 
        blank17_7, blank17_NE_3, \frame_begin[5]_net_1 , 
        \counter[5]_net_1 , blank17_6, blank17_NE_2, 
        \frame_begin[4]_net_1 , blank17_3, blank17_NE_1, blank17_2, 
        \counter[9]_net_1 , \frame_begin[9]_net_1 , awaitscheme7_2, 
        un1_data_sent_NE_13, un1_data_sent_NE_5, un1_data_sent_NE_4, 
        un1_data_sent_NE_11, un1_data_sent_NE_12, un1_data_sent_NE_3, 
        un1_data_sent_NE_2, un1_data_sent_NE_8, un1_data_sent_5, 
        un1_data_sent_4, un1_data_sent_NE_7, un1_data_sent_9, 
        un1_data_sent_8, un1_data_sent_NE_1, \data_sent[6]_net_1 , 
        \data_size[6]_net_1 , un1_data_sent_7, \data_sent[2]_net_1 , 
        \data_size[2]_net_1 , un1_data_sent_3, \data_sent[0]_net_1 , 
        \data_size[0]_net_1 , un1_data_sent_1, \data_sent[14]_net_1 , 
        \data_size[14]_net_1 , un1_data_sent_15, \data_sent[12]_net_1 , 
        \data_size[12]_net_1 , un1_data_sent_13, \data_sent[10]_net_1 , 
        \data_size[10]_net_1 , un1_data_sent_11, 
        awaitscheme_6_0_0_o2_0_0, N_248_i, \i[1]_net_1 , 
        awaitheartbeat_1_sqmuxa_1_0_o2_1, \counter[3]_net_1 , 
        awaitheartbeat_1_sqmuxa_1_0_o2_0, 
        data_size_1_sqmuxa_i_0_o2_4_2, \tick[7]_net_1 , 
        data_size_1_sqmuxa_i_0_o2_4_1, \tick[3]_net_1 , 
        data_size_1_sqmuxa_i_0_o2_4_0, \tick[9]_net_1 , 
        \tick[5]_net_1 , \counter[7]_net_1 , 
        un1_tick_0_sqmuxa_1_0_a2_4_1, un1_tick_0_sqmuxa_1_0_a2_4_0, 
        sending13_2, \data_len[5]_net_1 , \data_len[6]_net_1 , 
        sending13_1, \data_len[3]_net_1 , \data_len[4]_net_1 , 
        sending13_0, \data_len[7]_net_1 , \data_len[8]_net_1 , N_269, 
        N_403, N_513, N_283, N_265, N_325, N_158, N_405, N_408, N_16, 
        N_363, N_355, N_46, \un1_frame_begin[6] , N_55, N_411, N_410, 
        N_409, un1_start_1_sqmuxa_3, N_299, rd_0_sqmuxa, N_338, N_370, 
        \un1_frame_begin[5] , \un1_choice_2[5] , I4_un1_CO1, 
        \un1_choice_2[6] , \frame_begin[6]_net_1 , N147, 
        calculating_0_sqmuxa, un1_calculating_0_sqmuxa, rd_0_sqmuxa_1, 
        N_287, un1_tick_0_sqmuxa, N_304, N_256, N_379, N_358, N_380, 
        I_35_0, N_464, N_413, \tick_14[4] , \tick_14_0_0_0[4] , N_504, 
        N_244, N_340, N_457, N_456, N_432, N_14, N_66, 
        un1_resuming_0_sqmuxa_5, N_386, resuming_0_sqmuxa_2, N_320, 
        N_268, \un1_frame_begin[4] , \un1_choice_2[4] , N143, N_415, 
        N_52, N_414, N_50, N_48, N_875, N_297, un1_start_1_sqmuxa_7, 
        N_874, \i[0]_net_1 , N_474, ie, N_423, i_0_sqmuxa, N_251, 
        un1_start_1_sqmuxa_4, N_200, counting_0_sqmuxa, cnt_n2, cnt_c1, 
        cnt_n3, cnt_c2, resuming_0_sqmuxa, un1_start_1_sqmuxa, N_396, 
        N_395, un1_start_1_sqmuxa_1, counting_0_sqmuxa_1, N_395_1, 
        un1_start_1_sqmuxa_2, i_1_sqmuxa, flag_1_sqmuxa, 
        \tick_14_0_0_a3_2_2[4] , cnt_n1_0_tz, cnt_c0, cnt_n0_0_tz, 
        cnt_n1, cnt_n0, un1_tick_0_sqmuxa_1, un1_tick_0_sqmuxa_1_1_0, 
        I8_un1_CO1, N151, I6_un1_CO1, \un1_choice_2[3] , 
        \frame_begin_18[3] , N_63, \frame_begin_18[7] , 
        \frame_begin_18[8] , \div_counter_3[1] , I_5_0, 
        \div_counter_3[4] , I_12_1, \div_counter_3[5] , I_14_1, N_378, 
        \frame_begin[2]_net_1 , \memo[1]_net_1 , un1_ord_0, 
        \flag_14[6] , \flag[7]_net_1 , \randint_12[7] , 
        \randint[10]_net_1 , \randint_12[10] , \randint[13]_net_1 , 
        \randint_12[12] , \randint[15]_net_1 , \randint_12[14] , 
        \randint[17]_net_1 , \randint_12[15] , \randint[18]_net_1 , 
        \randint_12[17] , \randint[20]_net_1 , \randint_12[18] , 
        \randint[21]_net_1 , \randint_12[19] , \randint[22]_net_1 , 
        \randint_12[20] , \randint[23]_net_1 , \scheme_11[0] , 
        \scheme[6]_net_1 , \scheme_11[2] , \scheme[8]_net_1 , 
        \scheme_11[3] , \scheme[9]_net_1 , \scheme_11[6] , 
        \scheme[12]_net_1 , \scheme_11[9] , \scheme[15]_net_1 , 
        \scheme_11[10] , \scheme[16]_net_1 , \scheme_11[11] , 
        \scheme[17]_net_1 , \scheme_11[12] , \scheme[18]_net_1 , 
        \scheme_11[13] , \scheme[19]_net_1 , \scheme_11[14] , 
        \scheme[20]_net_1 , \scheme_11[15] , \scheme[21]_net_1 , 
        \scheme_11[16] , \scheme[22]_net_1 , \scheme_11[17] , 
        \scheme[23]_net_1 , \scheme_11[18] , \scheme[24]_net_1 , 
        \scheme_11[19] , \scheme[25]_net_1 , \scheme_11[20] , 
        \scheme[26]_net_1 , \scheme_11[21] , \scheme[27]_net_1 , 
        \scheme_11[22] , \scheme[28]_net_1 , \scheme_11[23] , 
        \scheme[29]_net_1 , \scheme_11[24] , \scheme[30]_net_1 , 
        \scheme_11[26] , \scheme[32]_net_1 , \scheme_11[27] , 
        \scheme[33]_net_1 , \scheme_11[28] , \scheme[34]_net_1 , 
        \scheme_11[29] , \scheme[35]_net_1 , \scheme_11[30] , 
        \scheme[36]_net_1 , \scheme_11[31] , \scheme[37]_net_1 , 
        \scheme_11[32] , \scheme[38]_net_1 , \scheme_11[33] , 
        \scheme[39]_net_1 , \scheme_11[34] , \scheme[40]_net_1 , 
        \scheme_11[35] , \scheme[41]_net_1 , \scheme_11[36] , 
        \scheme[42]_net_1 , \scheme_11[37] , \scheme[43]_net_1 , 
        \scheme_11[38] , \scheme[44]_net_1 , \scheme_11[39] , 
        \scheme[45]_net_1 , \scheme_11[40] , \scheme[46]_net_1 , 
        \scheme_11[41] , \scheme[47]_net_1 , \randint_12[4] , 
        \randint[7]_net_1 , \randint_12[5] , \randint[8]_net_1 , 
        \randint_12[11] , \randint[14]_net_1 , \randint_12[8] , 
        \randint[11]_net_1 , \data_size[1]_net_1 , 
        \data_sent[1]_net_1 , data_sent_e0, data_sent_1_sqmuxa_1, 
        \data_size[3]_net_1 , \data_sent[3]_net_1 , 
        \data_size[4]_net_1 , \data_sent[4]_net_1 , 
        \data_size[5]_net_1 , \data_sent[5]_net_1 , 
        \data_size[7]_net_1 , \data_sent[7]_net_1 , 
        \data_size[8]_net_1 , \data_sent[8]_net_1 , 
        \data_size[9]_net_1 , \data_sent[9]_net_1 , 
        \data_size[11]_net_1 , \data_sent[11]_net_1 , 
        \data_size[13]_net_1 , \data_sent[13]_net_1 , 
        \data_sent[15]_net_1 , \data_size[15]_net_1 , data_sent_n15, 
        data_sent_c13, \memo[0]_net_1 , data_sent_n14, data_sent_n13, 
        data_sent_c12, data_sent_n12, data_sent_c10, data_sent_n11, 
        data_sent_n10, data_sent_c8, data_sent_n9, data_sent_n8, 
        data_sent_c6, data_sent_n7, data_sent_n6, data_sent_c4, 
        data_sent_n5, data_sent_n4, data_sent_c2, data_sent_n3, 
        data_sent_n2, data_sent_n1, awaitheartbeat_RNO_net_1, i44, 
        N_508, \choice[0]_net_1 , \data_len_11[3] , \scheme[0]_net_1 , 
        \data_len_11[4] , \scheme[1]_net_1 , \data_len_11[5] , 
        \scheme[2]_net_1 , \data_len_11[6] , \scheme[3]_net_1 , 
        \data_len_11[7] , \scheme[4]_net_1 , N_393, N_434, 
        \data_len_11[8] , \scheme[5]_net_1 , N_458, N_487, N_149, 
        \counter_17[5] , I_34, un1_tick_2_sqmuxa_14, \counter_17[7] , 
        I_39, \counter_17[9] , I_38, N_239, N_344, N_345, N_346, N_348, 
        N_349, \flag_14[0] , \flag[1]_net_1 , \flag_14[7] , 
        \counter[0]_net_1 , \scheme_11[7] , \scheme[13]_net_1 , 
        \scheme_11[5] , \scheme[11]_net_1 , \scheme_11[4] , 
        \scheme[10]_net_1 , \frame_begin_18[9] , \counter_17[6] , I_36, 
        N_483, init_0_RNI7DURC2_net_1, \tick_14[2] , I_42_0, N_213, 
        \tick_14[9] , I_38_0, \tick_14[8] , I_40_0, \tick_14[7] , 
        I_39_0, \tick_14[6] , I_36_0, \tick_14[5] , I_34_0, 
        \tick_14[3] , I_33_0, \tick_14[1] , I_37_0, \tick_14[0] , 
        \DWACT_ADD_CI_0_partial_sum[0] , data_sent_1_sqmuxa_1_1, 
        awaitscheme_net_1, awaitscheme_6, N_67, N_328, N_336, 
        \id[2]_net_1 , N_278, un1_frame_begin_0_sqmuxa, N_444, N_315, 
        N_114, N_873, \counter_17[8] , I_40, \counter_17[4] , I_35, 
        \counter_17[3] , I_33, \counter_17[2] , I_42, \counter_17[1] , 
        I_37, \counter_17[0] , \DWACT_ADD_CI_0_partial_sum_0[0] , 
        \flag_14[2] , \flag[3]_net_1 , \flag_14[1] , \flag[2]_net_1 , 
        N_347, \scheme_11[25] , \scheme[31]_net_1 , \scheme_11[8] , 
        \scheme[14]_net_1 , un1_tick_2_sqmuxa_3, un1_start_1_sqmuxa_6, 
        un1_resuming_0_sqmuxa_3, N_526, un1_counting_0_sqmuxa, 
        un1_start_0_sqmuxa, N_495, \DWACT_ADD_CI_0_partial_sum_1[0] , 
        \randint[0]_net_1 , N_496, I_12_0, \randint[1]_net_1 , N_497, 
        I_14_0, \randint[2]_net_1 , \rd_13[0] , \rd_13[1] , \rd_13[2] , 
        \randint_12[21] , \randint_12[2] , \randint[5]_net_1 , 
        \randint_12[1] , \randint[4]_net_1 , \randint_12[0] , 
        \randint[3]_net_1 , \randint_12[23] , \randint_12[22] , 
        \randint_12[16] , \randint[19]_net_1 , \randint_12[13] , 
        \randint[16]_net_1 , \randint_12[9] , \randint[12]_net_1 , 
        \randint_12[6] , \randint[9]_net_1 , \randint_12[3] , 
        \randint[6]_net_1 , \flag_14[5] , \flag[6]_net_1 , 
        \scheme_11[1] , \scheme[7]_net_1 , \flag_14[4] , 
        \flag[5]_net_1 , \flag_14[3] , \flag[4]_net_1 , \id[0]_net_1 , 
        \id[1]_net_1 , I_4_0, I_7_0, I_9_0, 
        \DWACT_ADD_CI_0_g_array_1_1[0] , 
        \DWACT_ADD_CI_0_pog_array_0[0] , \DWACT_ADD_CI_0_TMP_1[0] , 
        \DWACT_ADD_CI_0_g_array_0_1[0] , 
        \DWACT_ADD_CI_0_partial_sum[2] , 
        \DWACT_ADD_CI_0_partial_sum[1] , N_2, N_4, 
        \DWACT_ADD_CI_0_pog_array_1_2[0] , 
        \DWACT_ADD_CI_0_pog_array_1_2_0[0] , GND, VCC;
    
    DFN1E1C0 \data_sent[12]  (.D(data_sent_n12), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[12]_net_1 ));
    DFN1 \cnt[0]  (.D(cnt_n0), .CLK(ref_signal_c), .Q(\cnt[0]_net_1 ));
    INV un3_div_counter_I_4 (.A(\div_counter[0]_net_1 ), .Y(I_4_0));
    DFN1P0 init_1 (.D(N_42), .CLK(ref_signal_c), .PRE(reset_c), .Q(
        init_1_net_1));
    OR2A \tick_RNIB7I34[4]  (.A(N_292), .B(N_274), .Y(
        id_1_sqmuxa_1_i_0_0));
    DFN1E1 \data_len[3]  (.D(\data_len_11[3] ), .CLK(ref_signal_c), .E(
        un1_frame_begin_0_sqmuxa), .Q(\data_len[3]_net_1 ));
    NOR3B past_RNISESB1 (.A(past_net_1), .B(reset_c), .C(N_264), .Y(
        un1_tick_2_sqmuxa_5_0_a2_1));
    XOR2 \data_sent_RNO[9]  (.A(data_sent_c8), .B(\data_sent[9]_net_1 )
        , .Y(data_sent_n9));
    NOR3B working_RNO_0 (.A(memo26), .B(N_477), .C(N_309), .Y(N_411));
    DFN1P0 init_0 (.D(N_42), .CLK(ref_signal_c), .PRE(reset_c), .Q(
        init_0_net_1));
    DFN1E0C0 \data_size[15]  (.D(\data_size[14]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[15]_net_1 ));
    NOR3B past_RNO (.A(N_263), .B(N_476), .C(N_304), .Y(
        un1_tick_0_sqmuxa));
    DFN1E1 \flag[1]  (.D(\flag_14[1] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_2), .Q(\flag[1]_net_1 ));
    NOR2B un1_counter_1_I_46 (.A(\DWACT_ADD_CI_0_g_array_1_0[0] ), .B(
        \counter[2]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12_0[0] ));
    DFN1E1 \flag[0]  (.D(\flag_14[0] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_2), .Q(\flag[0]_net_1 ));
    AND2 un1_counter_1_I_61 (.A(\DWACT_ADD_CI_0_pog_array_1_1_0[0] ), 
        .B(\DWACT_ADD_CI_0_pog_array_1_2[0] ), .Y(
        \DWACT_ADD_CI_0_pog_array_2_0[0] ));
    NOR2B un1_counter_1_I_47 (.A(\DWACT_ADD_CI_0_g_array_2_0[0] ), .B(
        \counter[4]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12_1_0[0] ));
    NOR3B init_RNI66M55 (.A(memo26), .B(N_480), .C(N_309), .Y(N_410));
    NOR3 init_0_RNISD4C5 (.A(init_0_net_1), .B(N_251), .C(N_291), .Y(
        N_483));
    MX2 \randint_RNO[12]  (.A(\randint[15]_net_1 ), .B(
        randgen_0_cur_rand[12]), .S(init_0_net_1), .Y(\randint_12[12] )
        );
    DFN1C0 \div_counter[4]  (.D(\div_counter_3[4] ), .CLK(ref_signal_c)
        , .CLR(reset_c), .Q(\div_counter[4]_net_1 ));
    NOR2B un1_counter_1_I_53 (.A(\DWACT_ADD_CI_0_g_array_2_0[0] ), .B(
        \DWACT_ADD_CI_0_pog_array_2_0[0] ), .Y(
        \DWACT_ADD_CI_0_g_array_3_0[0] ));
    MX2 \randint_RNO[20]  (.A(\randint[23]_net_1 ), .B(
        randgen_0_cur_rand[20]), .S(init_1_net_1), .Y(\randint_12[20] )
        );
    OR3 \data_size_RNIOB2P[4]  (.A(un1_data_sent_5), .B(
        un1_data_sent_4), .C(un1_data_sent_NE_7), .Y(
        un1_data_sent_NE_11));
    DFN1E1 \randint[0]  (.D(\randint_12[0] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[0]_net_1 ));
    NOR2B \data_sent_RNIL61N2[13]  (.A(data_sent_c12), .B(
        \data_sent[13]_net_1 ), .Y(data_sent_c13));
    AND2 un1_rd_1_I_5 (.A(\rd[1]_net_1 ), .B(rd_0_sqmuxa), .Y(
        \DWACT_ADD_CI_0_g_array_0_1[0] ));
    NOR2A \randint_RNO[5]  (.A(\randint[8]_net_1 ), .B(init_net_1), .Y(
        \randint_12[5] ));
    DFN1E1C0 \data_sent[13]  (.D(data_sent_n13), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[13]_net_1 ));
    AO13 \cnt_RNO_0[3]  (.A(cnt_c1), .B(\cnt[2]_net_1 ), .C(
        cnt_0_sqmuxa), .Y(cnt_c2));
    OR2 \cnt_RNIJJ7CD[0]  (.A(N_526), .B(\cnt[0]_net_1 ), .Y(cnt_c0));
    OR3 awaitbeacon_RNIKKG13 (.A(N_244), .B(N_457), .C(N_456), .Y(
        N_274));
    NOR3C \div_counter_RNIVPT42[1]  (.A(div_counter11_1), .B(
        div_counter11_0), .C(div_counter11_2), .Y(div_counter11));
    OR2 launch_RNIPLP4M (.A(N_444), .B(tick_2_sqmuxa), .Y(
        un1_tick_2_sqmuxa_2));
    OR3 \data_size_RNIK3G91[8]  (.A(un1_data_sent_9), .B(
        un1_data_sent_8), .C(un1_data_sent_NE_1), .Y(
        un1_data_sent_NE_8));
    DFN1E1 \randint[8]  (.D(\randint_12[8] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[8]_net_1 ));
    DFN1E1 \scheme[35]  (.D(\scheme_11[35] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[35]_net_1 ));
    DFN1E1 \i[0]  (.D(N_873), .CLK(ref_signal_c), .E(ie), .Q(
        \i[0]_net_1 ));
    XOR2 un1_tick_3_I_36 (.A(\tick[6]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_11[0] ), .Y(I_36_0));
    DFN1E1 resuming (.D(un1_resuming_0_sqmuxa_3), .CLK(ref_signal_c), 
        .E(un1_resuming_0_sqmuxa_5), .Q(resuming_net_1));
    DFN1E1 \randint[9]  (.D(\randint_12[9] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[9]_net_1 ));
    MX2 \randint_RNO[9]  (.A(\randint[12]_net_1 ), .B(
        randgen_0_cur_rand[9]), .S(init_net_1), .Y(\randint_12[9] ));
    DFN1E1 \randint[5]  (.D(\randint_12[5] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[5]_net_1 ));
    MX2 \scheme_RNO[11]  (.A(\scheme[17]_net_1 ), .B(
        demodulator_0_cur_scheme[11]), .S(init_1_net_1), .Y(
        \scheme_11[11] ));
    OR2A init_RNIHI39F (.A(N_284), .B(N_385), .Y(
        un1_frame_begin_0_sqmuxa));
    DFN1E1 \scheme[37]  (.D(\scheme_11[37] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[37]_net_1 ));
    MX2 \rd_RNO_0[1]  (.A(I_12_0), .B(\randint[1]_net_1 ), .S(
        resuming_0_sqmuxa_2), .Y(N_496));
    DFN1E0C0 \data_size[11]  (.D(\data_size[10]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[11]_net_1 ));
    XOR2 un1_counter_1_I_36 (.A(\counter[6]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_11_0[0] ), .Y(I_36));
    XOR2 \data_sent_RNO[11]  (.A(data_sent_c10), .B(
        \data_sent[11]_net_1 ), .Y(data_sent_n11));
    OR3 \tick_RNIP6CR7[4]  (.A(data_size_1_sqmuxa_i_0_0), .B(N_265), 
        .C(N_355), .Y(N_14));
    DFN1E1C0 \data_sent[15]  (.D(data_sent_n15), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[15]_net_1 ));
    OA1B \counter_RNIAQ0V1[3]  (.A(N_500), .B(N_501), .C(N_287), .Y(
        N_370));
    NOR3A blank_RNIG7CJ (.A(blank_net_1), .B(init_0_net_1), .C(
        launch_net_1), .Y(start_2_sqmuxa_0));
    OR2 past_RNINI471 (.A(un1_tick_0_sqmuxa_1_0_0_o2_1), .B(N_287), .Y(
        N_291));
    XOR2 un1_counter_1_I_37 (.A(\counter[1]_net_1 ), .B(
        \DWACT_ADD_CI_0_TMP_0[0] ), .Y(I_37));
    MX2 \scheme_RNO[37]  (.A(\scheme[43]_net_1 ), .B(
        demodulator_0_cur_scheme[37]), .S(init_2_net_1), .Y(
        \scheme_11[37] ));
    AND2 un1_rd_1_I_1 (.A(\rd[0]_net_1 ), .B(rd_0_sqmuxa), .Y(
        \DWACT_ADD_CI_0_TMP_1[0] ));
    DFN1E1 \randint[14]  (.D(\randint_12[14] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[14]_net_1 ));
    NOR3C \data_sent_RNI19IV1[10]  (.A(\data_sent[9]_net_1 ), .B(
        data_sent_c8), .C(\data_sent[10]_net_1 ), .Y(data_sent_c10));
    AO1A past_RNO_0 (.A(N_251), .B(un1_tick_0_sqmuxa_1_0_0_0_0), .C(
        un1_tick_0_sqmuxa_1_1_0), .Y(un1_tick_0_sqmuxa_1));
    XOR2 \frame_begin_RNI10J6[3]  (.A(\counter[3]_net_1 ), .B(
        \frame_begin[3]_net_1 ), .Y(blank17_3));
    AO1 awaitscheme_RNO (.A(N_340), .B(awaitscheme_net_1), .C(N_413), 
        .Y(awaitscheme_6));
    XOR2 un1_rd_1_I_14 (.A(\DWACT_ADD_CI_0_partial_sum[2] ), .B(
        \DWACT_ADD_CI_0_g_array_1_1[0] ), .Y(I_14_0));
    NOR3C \memo_RNIHDSK6[1]  (.A(div_counter11), .B(memo26), .C(N_274), 
        .Y(N_403));
    XOR2 un1_counter_1_I_38 (.A(\counter[9]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12_3_0[0] ), .Y(I_38));
    DFN1 \frame_begin[2]  (.D(N_52), .CLK(ref_signal_c), .Q(
        \frame_begin[2]_net_1 ));
    DFN1E0C0 \data_size[14]  (.D(\data_size[13]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[14]_net_1 ));
    MX2 \flag_RNO[1]  (.A(\flag[2]_net_1 ), .B(
        demodulator_0_cur_flag[1]), .S(init_1_net_1), .Y(\flag_14[1] ));
    OR3 calculating_RNICL2I6 (.A(N_265), .B(N_269), .C(
        tick_1_sqmuxa_2_i_i_o2_0), .Y(N_283));
    NOR2B \tick_RNO[6]  (.A(I_36_0), .B(N_213), .Y(\tick_14[6] ));
    MX2 \scheme_RNO[19]  (.A(\scheme[25]_net_1 ), .B(
        demodulator_0_cur_scheme[19]), .S(init_2_net_1), .Y(
        \scheme_11[19] ));
    OAI1 blank_RNO (.A(N_464), .B(un1_tick_2_sqmuxa_0), .C(N_314), .Y(
        un1_tick_2_sqmuxa_3));
    OR3 \frame_begin_RNIF9DR[5]  (.A(blank17_NE_0), .B(blank17_7), .C(
        blank17_NE_3), .Y(blank17_NE_6));
    DFN1 \cnt[3]  (.D(cnt_n3), .CLK(ref_signal_c), .Q(\cnt[3]_net_1 ));
    NOR2B un1_tick_3_I_44 (.A(\DWACT_ADD_CI_0_g_array_3[0] ), .B(
        \tick[8]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12_3[0] ));
    MX2 \scheme_RNO[2]  (.A(\scheme[8]_net_1 ), .B(
        demodulator_0_cur_scheme[2]), .S(init_0_net_1), .Y(
        \scheme_11[2] ));
    AO1D \data_size_RNI9ALB5[0]  (.A(un1_data_sent_NE_13), .B(
        un1_data_sent_NE_12), .C(sending13), .Y(N_312));
    DFN1E1 \scheme[18]  (.D(\scheme_11[18] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[18]_net_1 ));
    DFN1E0C0 \data_size[9]  (.D(\data_size[8]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[9]_net_1 ));
    OR3A past_RNI14341 (.A(past_net_1), .B(start_net_1), .C(N_264), .Y(
        un1_tick_0_sqmuxa_1_0_0_o2_1));
    OR2 launch_RNO_1 (.A(start_1_sqmuxa), .B(tick_2_sqmuxa), .Y(
        un1_start_1_sqmuxa_4_0));
    XO1 \frame_begin_RNIA86D[8]  (.A(\frame_begin[8]_net_1 ), .B(
        \counter[8]_net_1 ), .C(blank17_2), .Y(blank17_NE_1));
    OA1B init_RNIDF1B3 (.A(N_500), .B(N_501), .C(N_309), .Y(
        memo_0_sqmuxa_1_i_i_a3_0));
    DFN1E1 \scheme[28]  (.D(\scheme_11[28] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[28]_net_1 ));
    NOR3A \counter_RNIQLVT_0[5]  (.A(N_245), .B(
        awaitscheme_6_0_0_o2_4_0), .C(awaitscheme_6_0_0_o2_4_1), .Y(
        N_501));
    MX2 \scheme_RNO[18]  (.A(\scheme[24]_net_1 ), .B(
        demodulator_0_cur_scheme[18]), .S(init_2_net_1), .Y(
        \scheme_11[18] ));
    XA1B \frame_begin_RNO[8]  (.A(N151), .B(ADD_10x10_slow_I8_S_0), .C(
        N_63), .Y(\frame_begin_18[8] ));
    XO1 \data_size_RNI8HGC[0]  (.A(\data_sent[0]_net_1 ), .B(
        \data_size[0]_net_1 ), .C(un1_data_sent_1), .Y(
        un1_data_sent_NE_4));
    XOR2 \data_size_RNI3O86[8]  (.A(\data_size[8]_net_1 ), .B(
        \data_sent[8]_net_1 ), .Y(un1_data_sent_8));
    DFN1P0 init_2 (.D(N_42), .CLK(ref_signal_c), .PRE(reset_c), .Q(
        init_2_net_1));
    OR3A launch_RNIECIE4 (.A(launch_net_1), .B(init_0_net_1), .C(N_251)
        , .Y(N_269));
    AOI1B awaitbeacon_RNO (.A(awaitbeacon_0_i_a3_0), .B(N_477), .C(
        awaitbeacon_net_1), .Y(N_239));
    NOR2A \randint_RNO[2]  (.A(\randint[5]_net_1 ), .B(init_net_1), .Y(
        \randint_12[2] ));
    NOR2B \tick_RNO[3]  (.A(I_33_0), .B(N_213), .Y(\tick_14[3] ));
    DFN1 \tick[8]  (.D(\tick_14[8] ), .CLK(ref_signal_c), .Q(
        \tick[8]_net_1 ));
    DFN1E1 \scheme[14]  (.D(\scheme_11[14] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[14]_net_1 ));
    NOR2A counting_RNIFHV81 (.A(N_472), .B(counting_net_1), .Y(N_479));
    NOR2A \randint_RNO[1]  (.A(\randint[4]_net_1 ), .B(init_net_1), .Y(
        \randint_12[1] ));
    DFN1E1 counting (.D(start_1_sqmuxa), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_1), .Q(counting_net_1));
    OR2A start_RNI669OC2 (.A(N_336), .B(N_432), .Y(N_213));
    MX2 \scheme_RNO[30]  (.A(\scheme[36]_net_1 ), .B(
        demodulator_0_cur_scheme[30]), .S(init_2_net_1), .Y(
        \scheme_11[30] ));
    OA1B past_RNO_1 (.A(N_477), .B(N_480), .C(N_291), .Y(
        un1_tick_0_sqmuxa_1_0_0_0_0));
    NOR3A \flag_RNIF92A6[0]  (.A(N_487), .B(N_265), .C(N_269), .Y(
        resuming_0_sqmuxa));
    DFN1E0C0 \data_size[6]  (.D(\data_size[5]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[6]_net_1 ));
    AND2 sending_7_i_i_a3_1 (.A(N_884), .B(sending_7_i_i_a3_1_0_net_1), 
        .Y(N_407));
    DFN1E1 \scheme[24]  (.D(\scheme_11[24] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[24]_net_1 ));
    OR2 calculating_RNO_0 (.A(un1_calculating_0_sqmuxa_0_0_0), .B(
        rd_0_sqmuxa_1), .Y(un1_calculating_0_sqmuxa));
    MAJ3 un1_frame_begin_ADD_10x10_slow_I3_CO1 (.A(
        \frame_begin[3]_net_1 ), .B(\un1_choice_2[3] ), .C(I2_un1_CO1), 
        .Y(N143));
    DFN1E1 \choice[0]  (.D(\i[0]_net_1 ), .CLK(ref_signal_c), .E(
        rd_0_sqmuxa_1), .Q(\choice[0]_net_1 ));
    OR2 \tick_RNIDVP6[3]  (.A(\tick[8]_net_1 ), .B(\tick[3]_net_1 ), 
        .Y(data_size_1_sqmuxa_i_0_o2_4_1));
    DFN1E0 blank (.D(N_464), .CLK(ref_signal_c), .E(
        un1_tick_2_sqmuxa_3), .Q(blank_net_1));
    OR2A \i_RNIGDOOD[1]  (.A(N_259), .B(N_200), .Y(N_314));
    DFN1E0C0 \data_size[8]  (.D(\data_size[7]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[8]_net_1 ));
    XOR2 un1_rd_1_I_11 (.A(\rd[1]_net_1 ), .B(rd_0_sqmuxa), .Y(
        \DWACT_ADD_CI_0_partial_sum[1] ));
    NOR2 \tick_RNIIKKU[2]  (.A(N_278), .B(N_268), .Y(N_476));
    DFN1E1C0 working (.D(N_55), .CLK(ref_signal_c), .CLR(reset_c), .E(
        div_counter11), .Q(mac_0_working));
    DFN1E1 \scheme[8]  (.D(\scheme_11[8] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[8]_net_1 ));
    DFN1 \frame_begin[4]  (.D(N_50), .CLK(ref_signal_c), .Q(
        \frame_begin[4]_net_1 ));
    OR3 counting_RNIGTI2K_0 (.A(N_401), .B(start_1_sqmuxa), .C(N_400), 
        .Y(un1_start_1_sqmuxa_3));
    OR3A awaitbeacon_RNI7Q3F1 (.A(demodulator_0_ctg[1]), .B(
        awaitscheme_6_0_0_o2_0_0), .C(demodulator_0_ctg[0]), .Y(N_281));
    DFN1E1 \scheme[42]  (.D(N_344), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[42]_net_1 ));
    DFN1E1 \scheme[39]  (.D(\scheme_11[39] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[39]_net_1 ));
    NOR2B \div_counter_RNIPCVM[5]  (.A(\div_counter[5]_net_1 ), .B(
        \div_counter[4]_net_1 ), .Y(div_counter11_0));
    OR3 awaitscheme_RNO_2 (.A(awaitscheme_6_0_0_o2_4_0), .B(
        awaitscheme_6_0_0_o2_4_1), .C(N_281), .Y(
        awaitscheme_6_0_0_o2_0));
    MAJ3 un1_frame_begin_ADD_10x10_slow_I7_CO1 (.A(
        \frame_begin[7]_net_1 ), .B(I6_un1_CO1), .C(\un1_choice_2[7] ), 
        .Y(N151));
    NOR2A awaitscheme_RNIHRSV (.A(N_252), .B(demodulator_0_ctg[1]), .Y(
        N_457));
    DFN1E1C0 \data_sent[14]  (.D(data_sent_n14), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[14]_net_1 ));
    OR2A launch_RNO (.A(N_314), .B(start_1_sqmuxa), .Y(
        un1_start_1_sqmuxa_6));
    NOR3A counting_RNII2AM7 (.A(\un1_choice_2_0_a2_0[3] ), .B(N_281), 
        .C(N_269), .Y(N_474));
    OR3A \tick_RNINI121[0]  (.A(\tick[0]_net_1 ), .B(\tick[1]_net_1 ), 
        .C(N_288), .Y(N_325));
    DFN1E1 \flag[5]  (.D(\flag_14[5] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_2), .Q(\flag[5]_net_1 ));
    AO1 calculating_RNO_1 (.A(un1_calculating_0_sqmuxa_0_0_a3_0), .B(
        N_482), .C(start_1_sqmuxa), .Y(un1_calculating_0_sqmuxa_0_0_0));
    OR3 blank_RNIIHK14 (.A(N_465), .B(blank_net_1), .C(N_509), .Y(
        sending_7_i_i_o2_0_1));
    OR2A \counter_RNISP01[9]  (.A(\counter[9]_net_1 ), .B(
        \counter[7]_net_1 ), .Y(awaitscheme_6_0_0_o2_4_0));
    NOR2A \tick_RNIPS8H1[4]  (.A(\tick[4]_net_1 ), .B(N_265), .Y(N_458)
        );
    DFN1E1 \randint[4]  (.D(\randint_12[4] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[4]_net_1 ));
    XOR2 \data_size_RNIRF86[4]  (.A(\data_size[4]_net_1 ), .B(
        \data_sent[4]_net_1 ), .Y(un1_data_sent_4));
    DFN1E1 \flag[2]  (.D(\flag_14[2] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_2), .Q(\flag[2]_net_1 ));
    MX2 \rd_RNO_0[2]  (.A(I_14_0), .B(\randint[2]_net_1 ), .S(
        resuming_0_sqmuxa_2), .Y(N_497));
    MX2 \scheme_RNO[32]  (.A(\scheme[38]_net_1 ), .B(
        demodulator_0_cur_scheme[32]), .S(init_2_net_1), .Y(
        \scheme_11[32] ));
    OA1 counting_RNITRJO1 (.A(un1_resuming_0_sqmuxa_5_0_0_o2_0), .B(
        un1_resuming_0_sqmuxa_5_0_0_o2_1), .C(counting_net_1), .Y(
        \un1_choice_2_0_a2_0[3] ));
    NOR2A \tick_RNIUPVT1_0[4]  (.A(N_245), .B(N_292), .Y(N_509));
    DFN1E1C0 \data_sent[5]  (.D(data_sent_n5), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[5]_net_1 ));
    XOR2 \data_sent_RNO[5]  (.A(data_sent_c4), .B(\data_sent[5]_net_1 )
        , .Y(data_sent_n5));
    NOR2B \scheme_RNI2BHS7[5]  (.A(\scheme[5]_net_1 ), .B(N_474), .Y(
        \un1_choice_2[8] ));
    DFN1E1 \flag[7]  (.D(\flag_14[7] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_2), .Q(\flag[7]_net_1 ));
    XOR2 \data_sent_RNO[0]  (.A(\data_sent[0]_net_1 ), .B(
        data_sent_1_sqmuxa_1), .Y(data_sent_e0));
    MX2 \scheme_RNO[33]  (.A(\scheme[39]_net_1 ), .B(
        demodulator_0_cur_scheme[33]), .S(init_2_net_1), .Y(
        \scheme_11[33] ));
    DFN1 \frame_begin[9]  (.D(\frame_begin_18[9] ), .CLK(ref_signal_c), 
        .Q(\frame_begin[9]_net_1 ));
    OR3A \counter_RNIME13[3]  (.A(awaitscheme7_2), .B(
        awaitheartbeat_1_sqmuxa_1_0_o2_1), .C(
        awaitheartbeat_1_sqmuxa_1_0_o2_0), .Y(N_287));
    DFN1E1 \randint[22]  (.D(\randint_12[22] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[22]_net_1 ));
    NOR2A \data_len_RNO[6]  (.A(\scheme[3]_net_1 ), .B(
        demodulator_0_ctg[0]), .Y(\data_len_11[6] ));
    NOR2 \flag_RNIOPPAD[0]  (.A(resuming_0_sqmuxa), .B(cnt_0_sqmuxa), 
        .Y(N_526));
    NOR3B awaitbeacon_RNIRRET3 (.A(demodulator_0_ctg[0]), .B(
        demodulator_0_ctg[1]), .C(N_274), .Y(tick_2_sqmuxa_1));
    DFN1E0C0 \data_size[10]  (.D(\data_size[9]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[10]_net_1 ));
    AO1A init_RNIRL9JD (.A(N_249), .B(memo_0_sqmuxa_1_i_i_a3_0), .C(
        N_403), .Y(N_149));
    MX2 awaitscheme_RNIGQSV (.A(awaitheartbeat_net_1), .B(
        awaitscheme_net_1), .S(demodulator_0_ctg[0]), .Y(N_244));
    XOR2 \data_sent_RNO[3]  (.A(data_sent_c2), .B(\data_sent[3]_net_1 )
        , .Y(data_sent_n3));
    OR2 init_RNIP32F1 (.A(N_291), .B(init_net_1), .Y(N_309));
    NOR3A blank_RNIOUNL7 (.A(start_2_sqmuxa_0), .B(N_274), .C(N_251), 
        .Y(start_2_sqmuxa));
    DFN1E1 \scheme[2]  (.D(\scheme_11[2] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[2]_net_1 ));
    DFN1E1 \randint[1]  (.D(\randint_12[1] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[1]_net_1 ));
    DFN1E1 \flag[4]  (.D(\flag_14[4] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_2), .Q(\flag[4]_net_1 ));
    MX2 \scheme_RNO[36]  (.A(\scheme[42]_net_1 ), .B(
        demodulator_0_cur_scheme[36]), .S(init_2_net_1), .Y(
        \scheme_11[36] ));
    DFN1E1 \randint[19]  (.D(\randint_12[19] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[19]_net_1 ));
    NOR2A \tick_RNIUPVT1[0]  (.A(id_1_sqmuxa_1_i_0_a2_0), .B(N_288), 
        .Y(N_513));
    OR3 sending_RNO (.A(N_405), .B(sending_7_i_i_0), .C(N_408), .Y(
        N_158));
    AO1 \counter_RNO[7]  (.A(I_39), .B(un1_tick_2_sqmuxa_14), .C(N_505)
        , .Y(\counter_17[7] ));
    MX2 \randint_RNO[10]  (.A(\randint[13]_net_1 ), .B(
        randgen_0_cur_rand[10]), .S(init_0_net_1), .Y(\randint_12[10] )
        );
    DFN1E1 start (.D(start_0_sqmuxa), .CLK(ref_signal_c), .E(
        un1_start_0_sqmuxa), .Q(start_net_1));
    XA1C \i_RNO[3]  (.A(\i[3]_net_1 ), .B(N_315), .C(
        un1_start_1_sqmuxa_7), .Y(N_114));
    DFN1 \tick[3]  (.D(\tick_14[3] ), .CLK(ref_signal_c), .Q(
        \tick[3]_net_1 ));
    OR3 resuming_RNO_0 (.A(N_386), .B(un1_resuming_0_sqmuxa_5_0_0_0), 
        .C(resuming_0_sqmuxa_2), .Y(un1_resuming_0_sqmuxa_5));
    GND GND_i (.Y(GND));
    DFN1E1 \scheme[7]  (.D(\scheme_11[7] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[7]_net_1 ));
    OR2A start_RNIRDTK (.A(start_net_1), .B(N_264), .Y(N_276));
    DFN1E1 \scheme[32]  (.D(\scheme_11[32] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[32]_net_1 ));
    OR2A \i_RNO_0[3]  (.A(\i[2]_net_1 ), .B(N_297), .Y(N_315));
    OR2 \counter_RNIOL01[8]  (.A(\counter[4]_net_1 ), .B(
        \counter[8]_net_1 ), .Y(awaitheartbeat_1_sqmuxa_1_0_o2_0));
    NOR2B \counter_RNO[2]  (.A(I_42), .B(un1_tick_2_sqmuxa_14), .Y(
        \counter_17[2] ));
    NOR2B un1_counter_1_I_51 (.A(\DWACT_ADD_CI_0_g_array_2_0[0] ), .B(
        \DWACT_ADD_CI_0_pog_array_1_1_0[0] ), .Y(
        \DWACT_ADD_CI_0_g_array_11_0[0] ));
    NOR2 \data_len_RNI3OB7[3]  (.A(\data_len[3]_net_1 ), .B(
        \data_len[4]_net_1 ), .Y(sending13_1));
    DFN1E1 \scheme[0]  (.D(\scheme_11[0] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[0]_net_1 ));
    OR2A \memo_RNIK2R04[1]  (.A(reset_c), .B(N_249), .Y(N_251));
    XOR2 \data_size_RNIL986[1]  (.A(\data_size[1]_net_1 ), .B(
        \data_sent[1]_net_1 ), .Y(un1_data_sent_1));
    OR2 resuming_RNO_2 (.A(N_385), .B(N_371), .Y(
        un1_resuming_0_sqmuxa_5_0_0_0));
    OA1C \frame_begin_RNO[5]  (.A(N_284), .B(\un1_frame_begin[5] ), .C(
        \frame_begin_18_i_0_0[5] ), .Y(N_48));
    NOR2A sending_RNO_3 (.A(mac_0_sending), .B(init_net_1), .Y(
        sending_7_i_i_a3_0_0));
    OR2B \memo_RNITOBJ3[1]  (.A(memo26), .B(div_counter11), .Y(N_249));
    DFN1 \frame_begin[8]  (.D(\frame_begin_18[8] ), .CLK(ref_signal_c), 
        .Q(\frame_begin[8]_net_1 ));
    NOR2A sending_7_i_i_a3_1_0 (.A(memo26), .B(N_329), .Y(
        sending_7_i_i_a3_1_0_net_1));
    NOR2B un1_tick_3_I_52 (.A(\DWACT_ADD_CI_0_g_array_11[0] ), .B(
        \tick[6]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12_2[0] ));
    MAJ3 un1_frame_begin_ADD_10x10_slow_I5_CO1 (.A(
        \frame_begin[5]_net_1 ), .B(I4_un1_CO1), .C(\un1_choice_2[5] ), 
        .Y(N147));
    DFN1E1 \randint[23]  (.D(\randint_12[23] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[23]_net_1 ));
    XO1 \i_RNI4VHN[3]  (.A(\i[1]_net_1 ), .B(\choice[1]_net_1 ), .C(
        \i[3]_net_1 ), .Y(un1_resuming_0_sqmuxa_5_0_0_o2_0));
    DFN1E1C0 \data_sent[11]  (.D(data_sent_n11), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[11]_net_1 ));
    NOR2B \tick_RNINI121_0[4]  (.A(N_476), .B(\tick[4]_net_1 ), .Y(
        N_478));
    AND3 un3_div_counter_I_8 (.A(\div_counter[0]_net_1 ), .B(
        \div_counter[1]_net_1 ), .C(\div_counter[2]_net_1 ), .Y(N_4));
    NOR2B sending_RNO_0 (.A(mac_0_sending), .B(N_299), .Y(N_405));
    AND3 un3_div_counter_I_13 (.A(\DWACT_FINC_E[0] ), .B(
        \div_counter[3]_net_1 ), .C(\div_counter[4]_net_1 ), .Y(N_2));
    MX2 \scheme_RNO[34]  (.A(\scheme[40]_net_1 ), .B(
        demodulator_0_cur_scheme[34]), .S(init_2_net_1), .Y(
        \scheme_11[34] ));
    OR3 \tick_RNIKT7R[2]  (.A(\tick[4]_net_1 ), .B(N_268), .C(
        \tick[2]_net_1 ), .Y(N_288));
    MX2 \scheme_RNO[15]  (.A(\scheme[21]_net_1 ), .B(
        demodulator_0_cur_scheme[15]), .S(init_1_net_1), .Y(
        \scheme_11[15] ));
    OR2 calculating_RNIEN0F7 (.A(N_283), .B(N_259), .Y(N_284));
    DFN1 \counter[0]  (.D(\counter_17[0] ), .CLK(ref_signal_c), .Q(
        \counter[0]_net_1 ));
    MX2 \scheme_RNO[0]  (.A(\scheme[6]_net_1 ), .B(
        demodulator_0_cur_scheme[0]), .S(init_0_net_1), .Y(
        \scheme_11[0] ));
    XO1 \memo_RNIUUDE1[1]  (.A(demodulator_0_ord[1]), .B(
        \memo[1]_net_1 ), .C(un1_ord_0), .Y(memo26));
    MX2 \randint_RNO[19]  (.A(\randint[22]_net_1 ), .B(
        randgen_0_cur_rand[19]), .S(init_1_net_1), .Y(\randint_12[19] )
        );
    DFN1 \counter[3]  (.D(\counter_17[3] ), .CLK(ref_signal_c), .Q(
        \counter[3]_net_1 ));
    MX2 \randint_RNO[7]  (.A(\randint[10]_net_1 ), .B(
        randgen_0_cur_rand[7]), .S(init_net_1), .Y(\randint_12[7] ));
    OR3 init_1_RNI19TP4 (.A(init_1_net_1), .B(N_251), .C(N_276), .Y(
        N_304));
    XOR2 un1_frame_begin_ADD_10x10_slow_I7_S_0 (.A(
        \frame_begin[7]_net_1 ), .B(\un1_choice_2[7] ), .Y(
        ADD_10x10_slow_I7_S_0));
    NOR2B init_RNI3R2Q7 (.A(un1_resuming_0_sqmuxa_5_0_0_a3_1), .B(
        N_443), .Y(N_385));
    NOR2B counting_RNIPGUP5 (.A(N_481), .B(counting_net_1), .Y(N_401));
    OR2 choosing_RNO (.A(counting_0_sqmuxa_1), .B(un1_start_1_sqmuxa_5)
        , .Y(un1_counting_0_sqmuxa));
    NOR2A launch_RNI981C8 (.A(tick_2_sqmuxa_1), .B(N_269), .Y(
        tick_2_sqmuxa));
    OR2B \i_RNIVUEE[1]  (.A(\i[1]_net_1 ), .B(\i[0]_net_1 ), .Y(N_297));
    OAI1 head_RNO_3 (.A(\tick[1]_net_1 ), .B(\tick[0]_net_1 ), .C(
        \id[2]_net_1 ), .Y(N_328));
    AX1C \data_sent_RNO[4]  (.A(\data_sent[3]_net_1 ), .B(data_sent_c2)
        , .C(\data_sent[4]_net_1 ), .Y(data_sent_n4));
    AO1 datacmd_RNO (.A(N_509), .B(N_312), .C(N_338), .Y(N_67));
    DFN1E1C0 \data_sent[10]  (.D(data_sent_n10), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[10]_net_1 ));
    NOR2B un3_div_counter_I_11 (.A(\div_counter[3]_net_1 ), .B(
        \DWACT_FINC_E[0] ), .Y(N_3));
    DFN1E0C0 \id[2]  (.D(\id[1]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_16), .Q(\id[2]_net_1 ));
    MX2 \scheme_RNO[47]  (.A(\scheme[5]_net_1 ), .B(
        demodulator_0_cur_scheme[47]), .S(init_net_1), .Y(N_349));
    OR3 \tick_RNO[4]  (.A(N_380), .B(\tick_14_0_0_0[4] ), .C(N_379), 
        .Y(\tick_14[4] ));
    MX2 \randint_RNO[3]  (.A(\randint[6]_net_1 ), .B(
        randgen_0_cur_rand[3]), .S(init_net_1), .Y(\randint_12[3] ));
    NOR2A \randint_RNO[8]  (.A(\randint[11]_net_1 ), .B(init_net_1), 
        .Y(\randint_12[8] ));
    OR2A \memo_RNIIJUF4[1]  (.A(memo26), .B(N_274), .Y(N_299));
    NOR3A counting_RNINDRS5 (.A(counting_net_1), .B(N_265), .C(N_269), 
        .Y(counting_0_sqmuxa));
    DFN1E1 \data_len[4]  (.D(\data_len_11[4] ), .CLK(ref_signal_c), .E(
        un1_frame_begin_0_sqmuxa), .Q(\data_len[4]_net_1 ));
    DFN1E1C0 \memo[0]  (.D(demodulator_0_ord[0]), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(N_149), .Q(\memo[0]_net_1 ));
    XA1C \cnt_RNO[1]  (.A(cnt_n1_0_tz), .B(cnt_0_sqmuxa), .C(
        un1_start_1_sqmuxa_5), .Y(cnt_n1));
    MX2 \randint_RNO[15]  (.A(\randint[18]_net_1 ), .B(
        randgen_0_cur_rand[15]), .S(init_0_net_1), .Y(\randint_12[15] )
        );
    NOR2A init_RNINECV (.A(un1_start_1_sqmuxa_1_0_0_a3_0), .B(
        init_net_1), .Y(un1_resuming_0_sqmuxa_5_0_0_a3_1));
    NOR3A launch_RNIHI9O5 (.A(launch_net_1), .B(N_251), .C(N_265), .Y(
        N_482));
    XA1C \i_RNO[2]  (.A(\i[2]_net_1 ), .B(N_297), .C(
        un1_start_1_sqmuxa_7), .Y(N_875));
    DFN1E1C0 \data_sent[8]  (.D(data_sent_n8), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[8]_net_1 ));
    DFN1E1 \randint[18]  (.D(\randint_12[18] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[18]_net_1 ));
    AND2 un1_counter_1_I_59 (.A(\counter[2]_net_1 ), .B(
        \counter[3]_net_1 ), .Y(\DWACT_ADD_CI_0_pog_array_1_0[0] ));
    MX2 \flag_RNO[0]  (.A(\flag[1]_net_1 ), .B(
        demodulator_0_cur_flag[0]), .S(init_1_net_1), .Y(\flag_14[0] ));
    OR3A \tick_RNI1JOFC[0]  (.A(N_363), .B(id_1_sqmuxa_1_i_0_0), .C(
        N_355), .Y(N_16));
    NOR2A \cnt_RNIOLR2[0]  (.A(\cnt[0]_net_1 ), .B(\cnt[2]_net_1 ), .Y(
        resuming_0_sqmuxa_2_0_a2_0_a3_1));
    OA1B awaitscheme_RNI03F01 (.A(demodulator_0_ctg[0]), .B(
        awaitscheme_net_1), .C(demodulator_0_ctg[1]), .Y(N_504));
    DFN1E1 \scheme[44]  (.D(N_346), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[44]_net_1 ));
    DFN1 \counter[7]  (.D(\counter_17[7] ), .CLK(ref_signal_c), .Q(
        \counter[7]_net_1 ));
    OR2A init_1_RNIPCS683 (.A(init_0_RNI7DURC2_net_1), .B(
        un1_tick_2_sqmuxa_5), .Y(un1_tick_2_sqmuxa_14));
    NOR2 data_sent_1_sqmuxa_1_0_a2_0_a2 (.A(N_312), .B(N_354), .Y(
        N_884));
    NOR2A counting_RNIPFPP6 (.A(counting_0_sqmuxa), .B(N_259), .Y(
        counting_0_sqmuxa_1));
    AX1C \data_sent_RNO[15]  (.A(\data_sent[14]_net_1 ), .B(
        data_sent_c13), .C(\data_sent[15]_net_1 ), .Y(data_sent_n15));
    AO1 awaitheartbeat_RNO (.A(N_410), .B(div_counter11), .C(
        awaitheartbeat_net_1), .Y(awaitheartbeat_RNO_net_1));
    NOR3C launch_RNILTEN (.A(counting_net_1), .B(launch_net_1), .C(
        reset_c), .Y(un1_start_1_sqmuxa_1_0_0_a3_0));
    XOR2 un1_tick_3_I_37 (.A(\tick[1]_net_1 ), .B(
        \DWACT_ADD_CI_0_TMP[0] ), .Y(I_37_0));
    NOR2 start_RNILKR012 (.A(N_274), .B(N_320), .Y(N_336));
    NOR2B un1_counter_1_I_52 (.A(\DWACT_ADD_CI_0_g_array_11_0[0] ), .B(
        \counter[6]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12_2_0[0] ));
    DFN1E1 \randint[2]  (.D(\randint_12[2] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[2]_net_1 ));
    DFN1E1 \choice[2]  (.D(\i[2]_net_1 ), .CLK(ref_signal_c), .E(
        rd_0_sqmuxa_1), .Q(\choice[2]_net_1 ));
    DFN1 \rd[2]  (.D(\rd_13[2] ), .CLK(ref_signal_c), .Q(\rd[2]_net_1 )
        );
    MX2 \scheme_RNO[27]  (.A(\scheme[33]_net_1 ), .B(
        demodulator_0_cur_scheme[27]), .S(init_2_net_1), .Y(
        \scheme_11[27] ));
    DFN1E1 \flag[6]  (.D(\flag_14[6] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_2), .Q(\flag[6]_net_1 ));
    NOR3C choosing_RNI8VH77 (.A(N_259), .B(N_395_1), .C(N_482), .Y(
        N_395));
    MX2 \scheme_RNO[9]  (.A(\scheme[15]_net_1 ), .B(
        demodulator_0_cur_scheme[9]), .S(init_0_net_1), .Y(
        \scheme_11[9] ));
    DFN1E1 \scheme[11]  (.D(\scheme_11[11] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[11]_net_1 ));
    NOR2 head_RNO (.A(head_13_0_i_0), .B(N_338), .Y(N_66));
    AO1D \frame_begin_RNO_0[6]  (.A(\choice[2]_net_1 ), .B(N_284), .C(
        N_505), .Y(\frame_begin_18_i_0_0[6] ));
    DFN1E1 \i[1]  (.D(N_874), .CLK(ref_signal_c), .E(ie), .Q(
        \i[1]_net_1 ));
    DFN1C0 \div_counter[3]  (.D(I_9_0), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\div_counter[3]_net_1 ));
    OA1 \tick_RNO_1[4]  (.A(\tick_14_0_0_a3_2_2[4] ), .B(N_320), .C(
        I_35_0), .Y(\tick_14_0_0_0[4] ));
    DFN1E1C0 \data_sent[4]  (.D(data_sent_n4), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[4]_net_1 ));
    DFN1E1 \scheme[21]  (.D(\scheme_11[21] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[21]_net_1 ));
    DFN1E0C0 \id[1]  (.D(\id[0]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_16), .Q(\id[1]_net_1 ));
    DFN1E0C0 \data_size[12]  (.D(\data_size[11]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[12]_net_1 ));
    MX2 \scheme_RNO[40]  (.A(\scheme[46]_net_1 ), .B(
        demodulator_0_cur_scheme[40]), .S(init_2_net_1), .Y(
        \scheme_11[40] ));
    NOR3A \cnt_RNIIDN5[3]  (.A(resuming_0_sqmuxa_2_0_a2_0_a3_1), .B(
        \cnt[1]_net_1 ), .C(\cnt[3]_net_1 ), .Y(
        resuming_0_sqmuxa_2_0_a2_0_a3_2));
    OR2 calculating_RNIAAKL (.A(calculating_net_1), .B(N_277), .Y(
        tick_1_sqmuxa_2_i_i_o2_0));
    XOR3 un1_frame_begin_ADD_10x10_slow_I4_S (.A(\un1_choice_2[4] ), 
        .B(\frame_begin[4]_net_1 ), .C(N143), .Y(\un1_frame_begin[4] ));
    DFN1 \tick[4]  (.D(\tick_14[4] ), .CLK(ref_signal_c), .Q(
        \tick[4]_net_1 ));
    MX2 \scheme_RNO[8]  (.A(\scheme[14]_net_1 ), .B(
        demodulator_0_cur_scheme[8]), .S(init_0_net_1), .Y(
        \scheme_11[8] ));
    NOR3 \frame_begin_RNO[2]  (.A(N_414), .B(N_505), .C(N_415), .Y(
        N_52));
    AND2 un1_tick_3_I_60 (.A(\tick[4]_net_1 ), .B(\tick[5]_net_1 ), .Y(
        \DWACT_ADD_CI_0_pog_array_1_1[0] ));
    NOR2B un1_tick_3_I_51 (.A(\DWACT_ADD_CI_0_g_array_2[0] ), .B(
        \DWACT_ADD_CI_0_pog_array_1_1[0] ), .Y(
        \DWACT_ADD_CI_0_g_array_11[0] ));
    DFN1E1 \scheme[38]  (.D(\scheme_11[38] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[38]_net_1 ));
    NOR2 \counter_RNIDA01[0]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(awaitscheme7_2));
    MX2 \scheme_RNO[6]  (.A(\scheme[12]_net_1 ), .B(
        demodulator_0_cur_scheme[6]), .S(init_0_net_1), .Y(
        \scheme_11[6] ));
    DFN1E1 \randint[20]  (.D(\randint_12[20] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[20]_net_1 ));
    DFN1E1C0 \data_sent[2]  (.D(data_sent_n2), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[2]_net_1 ));
    DFN1E1 \choice[1]  (.D(\i[1]_net_1 ), .CLK(ref_signal_c), .E(
        rd_0_sqmuxa_1), .Q(\choice[1]_net_1 ));
    NOR3B \tick_RNO_3[4]  (.A(N_292), .B(\tick_14_0_0_a3_2_2_0[4] ), 
        .C(N_304), .Y(\tick_14_0_0_a3_2_2[4] ));
    MX2A head_RNO_1 (.A(N_328), .B(\data_size[15]_net_1 ), .S(N_288), 
        .Y(N_361));
    OR2 \counter_RNIHE01[3]  (.A(\counter[2]_net_1 ), .B(
        \counter[3]_net_1 ), .Y(awaitheartbeat_1_sqmuxa_1_0_o2_1));
    AO1 \tick_RNISJVR3[0]  (.A(N_325), .B(N_245), .C(N_513), .Y(N_363));
    OR2 \tick_RNIF1Q6[7]  (.A(\tick[7]_net_1 ), .B(\tick[6]_net_1 ), 
        .Y(data_size_1_sqmuxa_i_0_o2_4_2));
    XOR2 \data_size_RNI5Q86[9]  (.A(\data_size[9]_net_1 ), .B(
        \data_sent[9]_net_1 ), .Y(un1_data_sent_9));
    OR3 counting_RNIGTI2K (.A(N_401), .B(start_1_sqmuxa), .C(N_400), 
        .Y(un1_start_1_sqmuxa_3_0));
    MX2 \scheme_RNO[31]  (.A(\scheme[37]_net_1 ), .B(
        demodulator_0_cur_scheme[31]), .S(init_2_net_1), .Y(
        \scheme_11[31] ));
    NOR2 awaitbeacon_RNO_0 (.A(N_309), .B(N_249), .Y(
        awaitbeacon_0_i_a3_0));
    DFN1P0 awaitbeacon (.D(N_239), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(awaitbeacon_net_1));
    NOR3A init_0_RNI8FU3A (.A(un1_tick_2_sqmuxa_5_0_a2_3), .B(N_370), 
        .C(N_299), .Y(N_154));
    NOR3B awaitscheme_RNO_1 (.A(memo26), .B(awaitscheme_6_0_0_a3_0_0), 
        .C(N_309), .Y(N_413));
    DFN1E1 \scheme[16]  (.D(\scheme_11[16] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[16]_net_1 ));
    OR2 \i_RNI22US[1]  (.A(un1_resuming_0_sqmuxa_3_0_0_o3_0), .B(N_256)
        , .Y(N_259));
    DFN1E1 \scheme[34]  (.D(\scheme_11[34] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[34]_net_1 ));
    MX2 \flag_RNO[6]  (.A(\flag[7]_net_1 ), .B(
        demodulator_0_cur_flag[6]), .S(init_1_net_1), .Y(\flag_14[6] ));
    NOR2B \counter_RNIOL01[5]  (.A(\counter[5]_net_1 ), .B(
        \counter[7]_net_1 ), .Y(un1_tick_0_sqmuxa_1_0_a2_4_1));
    MX2 \flag_RNO[2]  (.A(\flag[3]_net_1 ), .B(
        demodulator_0_cur_flag[2]), .S(init_1_net_1), .Y(\flag_14[2] ));
    XOR2 \data_sent_RNO[7]  (.A(data_sent_c6), .B(\data_sent[7]_net_1 )
        , .Y(data_sent_n7));
    NOR2A \div_counter_RNO[1]  (.A(I_5_0), .B(div_counter11), .Y(
        \div_counter_3[1] ));
    NOR2B un1_tick_3_I_55 (.A(\DWACT_ADD_CI_0_g_array_1[0] ), .B(
        \DWACT_ADD_CI_0_pog_array_1[0] ), .Y(
        \DWACT_ADD_CI_0_g_array_2[0] ));
    XNOR2 \cnt_RNO_0[0]  (.A(resuming_0_sqmuxa), .B(\cnt[0]_net_1 ), 
        .Y(cnt_n0_0_tz));
    NOR3A init_0_RNIPFG67 (.A(init_0_net_1), .B(N_274), .C(N_251), .Y(
        start_1_sqmuxa));
    DFN1E1 \scheme[26]  (.D(\scheme_11[26] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[26]_net_1 ));
    DFN1 \rd[1]  (.D(\rd_13[1] ), .CLK(ref_signal_c), .Q(\rd[1]_net_1 )
        );
    MX2 \scheme_RNO[20]  (.A(\scheme[26]_net_1 ), .B(
        demodulator_0_cur_scheme[20]), .S(init_2_net_1), .Y(
        \scheme_11[20] ));
    NOR2B un1_counter_1_I_56 (.A(\DWACT_ADD_CI_0_TMP_0[0] ), .B(
        \counter[1]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_1_0[0] ));
    XOR2 \data_size_RNIN9FE[11]  (.A(\data_size[11]_net_1 ), .B(
        \data_sent[11]_net_1 ), .Y(un1_data_sent_11));
    MX2 \scheme_RNO[42]  (.A(\scheme[0]_net_1 ), .B(
        demodulator_0_cur_scheme[42]), .S(init_net_1), .Y(N_344));
    DFN1E1 \i[3]  (.D(N_114), .CLK(ref_signal_c), .E(ie), .Q(
        \i[3]_net_1 ));
    AO1 counting_RNICF19E (.A(N_479), .B(N_481), .C(start_1_sqmuxa), 
        .Y(un1_start_1_sqmuxa_7_0_1_0));
    DFN1E0C0 \data_size[13]  (.D(\data_size[12]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[13]_net_1 ));
    MX2 \scheme_RNO[43]  (.A(\scheme[1]_net_1 ), .B(
        demodulator_0_cur_scheme[43]), .S(init_net_1), .Y(N_345));
    MX2 \scheme_RNO[4]  (.A(\scheme[10]_net_1 ), .B(
        demodulator_0_cur_scheme[4]), .S(init_0_net_1), .Y(
        \scheme_11[4] ));
    OR3 init_0_RNIVVVJK (.A(N_396), .B(start_1_sqmuxa), .C(N_395), .Y(
        un1_start_1_sqmuxa));
    NOR2A \tick_RNO_6[4]  (.A(demodulator_0_ctg[1]), .B(N_244), .Y(
        N_449));
    NOR3B \tick_RNO_0[4]  (.A(N_354), .B(I_35_0), .C(N_464), .Y(N_380));
    XOR2 \data_size_RNI1M86[7]  (.A(\data_size[7]_net_1 ), .B(
        \data_sent[7]_net_1 ), .Y(un1_data_sent_7));
    NOR3A sending_RNO_2 (.A(sending_7_i_i_a3_2_0), .B(N_299), .C(
        sending_7_i_i_o2_0_1), .Y(N_408));
    OR2 init_0_RNIQ6AMD (.A(resuming_0_sqmuxa_2), .B(start_1_sqmuxa), 
        .Y(un1_start_1_sqmuxa_5));
    DFN1 \tick[5]  (.D(\tick_14[5] ), .CLK(ref_signal_c), .Q(
        \tick[5]_net_1 ));
    MX2 \scheme_RNO[39]  (.A(\scheme[45]_net_1 ), .B(
        demodulator_0_cur_scheme[39]), .S(init_2_net_1), .Y(
        \scheme_11[39] ));
    DFN1E1 \randint[12]  (.D(\randint_12[12] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[12]_net_1 ));
    NOR2A \tick_RNIUPVT1[4]  (.A(N_478), .B(N_245), .Y(N_465));
    AND2 un1_counter_1_I_58 (.A(\counter[6]_net_1 ), .B(
        \counter[7]_net_1 ), .Y(\DWACT_ADD_CI_0_pog_array_1_2[0] ));
    DFN1E1 \scheme[9]  (.D(\scheme_11[9] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[9]_net_1 ));
    DFN1P0 init (.D(N_42), .CLK(ref_signal_c), .PRE(reset_c), .Q(
        init_net_1));
    NOR3A launch_RNI4EHP5 (.A(launch_net_1), .B(N_251), .C(N_281), .Y(
        N_481));
    NOR2B \choice_RNI5KOF7[0]  (.A(N_508), .B(\choice[0]_net_1 ), .Y(
        N_378));
    MX2 \scheme_RNO[46]  (.A(\scheme[4]_net_1 ), .B(
        demodulator_0_cur_scheme[46]), .S(init_net_1), .Y(N_348));
    AX1C \data_sent_RNO[10]  (.A(\data_sent[9]_net_1 ), .B(
        data_sent_c8), .C(\data_sent[10]_net_1 ), .Y(data_sent_n10));
    XOR2 un1_counter_1_I_35 (.A(\counter[4]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_2_0[0] ), .Y(I_35));
    OR2A init_0_RNIHI2BE (.A(N_284), .B(N_505), .Y(N_63));
    AO1 \scheme_RNI3R9CF[0]  (.A(\scheme[0]_net_1 ), .B(N_474), .C(
        N_393), .Y(\un1_choice_2[3] ));
    MX2 \scheme_RNO[38]  (.A(\scheme[44]_net_1 ), .B(
        demodulator_0_cur_scheme[38]), .S(init_2_net_1), .Y(
        \scheme_11[38] ));
    DFN1E1 \scheme[4]  (.D(\scheme_11[4] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[4]_net_1 ));
    NOR3 \tick_RNISHRJ8[4]  (.A(N_354), .B(N_312), .C(N_292), .Y(
        data_sent_1_sqmuxa_1_1));
    OR2 counting_RNO (.A(un1_start_1_sqmuxa_1_0_0_0), .B(
        counting_0_sqmuxa_1), .Y(un1_start_1_sqmuxa_1));
    DFN1E1 \scheme[13]  (.D(\scheme_11[13] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[13]_net_1 ));
    MX2 \scheme_RNO[22]  (.A(\scheme[28]_net_1 ), .B(
        demodulator_0_cur_scheme[22]), .S(init_2_net_1), .Y(
        \scheme_11[22] ));
    DFN1C0 \div_counter[5]  (.D(\div_counter_3[5] ), .CLK(ref_signal_c)
        , .CLR(reset_c), .Q(\div_counter[5]_net_1 ));
    DFN1E0 datacmd (.D(data_sent_1_sqmuxa_1_1), .CLK(ref_signal_c), .E(
        N_67), .Q(mac_0_datacmd));
    DFN1 \counter[2]  (.D(\counter_17[2] ), .CLK(ref_signal_c), .Q(
        \counter[2]_net_1 ));
    XOR2 un3_div_counter_I_5 (.A(\div_counter[0]_net_1 ), .B(
        \div_counter[1]_net_1 ), .Y(I_5_0));
    XOR3 un1_frame_begin_ADD_10x10_slow_I6_S (.A(\un1_choice_2[6] ), 
        .B(\frame_begin[6]_net_1 ), .C(N147), .Y(\un1_frame_begin[6] ));
    MX2 \scheme_RNO[23]  (.A(\scheme[29]_net_1 ), .B(
        demodulator_0_cur_scheme[23]), .S(init_2_net_1), .Y(
        \scheme_11[23] ));
    NOR2A \div_counter_RNO[4]  (.A(I_12_1), .B(div_counter11), .Y(
        \div_counter_3[4] ));
    DFN1E1C0 \data_sent[3]  (.D(data_sent_n3), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[3]_net_1 ));
    DFN1E0C0 \data_size[7]  (.D(\data_size[6]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[7]_net_1 ));
    DFN1E1 \scheme[23]  (.D(\scheme_11[23] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[23]_net_1 ));
    XOR2 \data_size_RNIPD86[3]  (.A(\data_size[3]_net_1 ), .B(
        \data_sent[3]_net_1 ), .Y(un1_data_sent_3));
    XOR2 \frame_begin_RNI76J6[6]  (.A(\counter[6]_net_1 ), .B(
        \frame_begin[6]_net_1 ), .Y(blank17_6));
    DFN1 \counter[6]  (.D(\counter_17[6] ), .CLK(ref_signal_c), .Q(
        \counter[6]_net_1 ));
    NOR2 \data_len_RNIB0C7[7]  (.A(\data_len[7]_net_1 ), .B(
        \data_len[8]_net_1 ), .Y(sending13_0));
    AO1 un1_rd_1_I_15 (.A(\DWACT_ADD_CI_0_pog_array_0[0] ), .B(
        \DWACT_ADD_CI_0_TMP_1[0] ), .C(\DWACT_ADD_CI_0_g_array_0_1[0] )
        , .Y(\DWACT_ADD_CI_0_g_array_1_1[0] ));
    NOR3A calculating_RNIQAIS (.A(calculating_net_1), .B(N_277), .C(
        \flag[0]_net_1 ), .Y(rd_0_sqmuxa_0));
    NOR2B un1_tick_3_I_46 (.A(\DWACT_ADD_CI_0_g_array_1[0] ), .B(
        \tick[2]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12[0] ));
    XOR2 un3_div_counter_I_12 (.A(N_3), .B(\div_counter[4]_net_1 ), .Y(
        I_12_1));
    OA1C working_RNO_1 (.A(init_1_net_1), .B(N_299), .C(mac_0_working), 
        .Y(N_409));
    XOR2 un3_div_counter_I_14 (.A(N_2), .B(\div_counter[5]_net_1 ), .Y(
        I_14_1));
    MX2 \flag_RNO[3]  (.A(\flag[4]_net_1 ), .B(
        demodulator_0_cur_flag[3]), .S(init_1_net_1), .Y(\flag_14[3] ));
    XO1 \data_size_RNIGPGC[2]  (.A(\data_sent[2]_net_1 ), .B(
        \data_size[2]_net_1 ), .C(un1_data_sent_3), .Y(
        un1_data_sent_NE_5));
    XOR2 un1_rd_1_I_10 (.A(\rd[2]_net_1 ), .B(rd_0_sqmuxa), .Y(
        \DWACT_ADD_CI_0_partial_sum[2] ));
    DFN1E1 \randint[13]  (.D(\randint_12[13] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[13]_net_1 ));
    DFN1E1 \scheme[10]  (.D(\scheme_11[10] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[10]_net_1 ));
    NOR2A blank_RNIDHGDL (.A(blank_net_1), .B(N_464), .Y(N_461));
    AO1 \scheme_RNI5T9CF[1]  (.A(\scheme[1]_net_1 ), .B(N_474), .C(
        N_434), .Y(\un1_choice_2[4] ));
    MX2 \scheme_RNO[26]  (.A(\scheme[32]_net_1 ), .B(
        demodulator_0_cur_scheme[26]), .S(init_2_net_1), .Y(
        \scheme_11[26] ));
    DFN1E1 \i[2]  (.D(N_875), .CLK(ref_signal_c), .E(ie), .Q(
        \i[2]_net_1 ));
    MX2 \scheme_RNO[44]  (.A(\scheme[2]_net_1 ), .B(
        demodulator_0_cur_scheme[44]), .S(init_net_1), .Y(N_346));
    NOR3C \data_len_RNILK3M[3]  (.A(sending13_1), .B(sending13_0), .C(
        sending13_2), .Y(sending13));
    DFN1E0C0 \data_size[5]  (.D(\data_size[4]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[5]_net_1 ));
    DFN1E1 \scheme[20]  (.D(\scheme_11[20] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[20]_net_1 ));
    AO1A init_0_RNI9PRBH (.A(N_251), .B(un1_start_0_sqmuxa_0_0_a3_1), 
        .C(start_1_sqmuxa), .Y(un1_tick_0_sqmuxa_1_1_0));
    NOR2B \counter_RNO[1]  (.A(I_37), .B(un1_tick_2_sqmuxa_14), .Y(
        \counter_17[1] ));
    XOR2 un1_tick_3_I_35 (.A(\tick[4]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_2[0] ), .Y(I_35_0));
    DFN1 \frame_begin[3]  (.D(\frame_begin_18[3] ), .CLK(ref_signal_c), 
        .Q(\frame_begin[3]_net_1 ));
    OR2A data_size_1_sqmuxa_i_0_o2 (.A(demodulator_0_ctg[0]), .B(
        demodulator_0_ctg[1]), .Y(N_245));
    OR3 init_0_RNIDOVKL (.A(i_1_sqmuxa), .B(start_1_sqmuxa), .C(
        flag_1_sqmuxa), .Y(un1_start_1_sqmuxa_2));
    OR3 \tick_RNINI121[4]  (.A(\tick[4]_net_1 ), .B(N_268), .C(N_278), 
        .Y(N_292));
    NOR3C \data_sent_RNIOR6F2[12]  (.A(\data_sent[11]_net_1 ), .B(
        data_sent_c10), .C(\data_sent[12]_net_1 ), .Y(data_sent_c12));
    NOR3A \tick_RNO_2[4]  (.A(N_358), .B(N_304), .C(N_265), .Y(N_379));
    OR2 init_1_RNILTDR7 (.A(N_304), .B(N_274), .Y(N_338));
    MX2 \randint_RNO[21]  (.A(\randint[0]_net_1 ), .B(
        randgen_0_cur_rand[21]), .S(init_1_net_1), .Y(\randint_12[21] )
        );
    MX2 \flag_RNO[4]  (.A(\flag[5]_net_1 ), .B(
        demodulator_0_cur_flag[4]), .S(init_1_net_1), .Y(\flag_14[4] ));
    NOR3A resuming_RNI2MN96 (.A(tick_1_sqmuxa_3_i_i_a3_0), .B(N_281), 
        .C(N_269), .Y(N_371));
    NOR2A \i_RNICCMQ6[3]  (.A(un1_resuming_0_sqmuxa_5_0_0_a2_0), .B(
        N_249), .Y(N_443));
    NOR2B \scheme_RNI09HS7[3]  (.A(\scheme[3]_net_1 ), .B(N_474), .Y(
        \un1_choice_2[6] ));
    XA1A \frame_begin_RNO_0[2]  (.A(\frame_begin[2]_net_1 ), .B(N_378), 
        .C(N_284), .Y(N_414));
    NOR2B \counter_RNO[3]  (.A(I_33), .B(un1_tick_2_sqmuxa_14), .Y(
        \counter_17[3] ));
    MX2 \rd_RNO_0[0]  (.A(\DWACT_ADD_CI_0_partial_sum_1[0] ), .B(
        \randint[0]_net_1 ), .S(resuming_0_sqmuxa_2), .Y(N_495));
    XA1B \frame_begin_RNO[3]  (.A(\un1_choice_2[3] ), .B(
        ADD_10x10_slow_I3_S_0), .C(N_63), .Y(\frame_begin_18[3] ));
    DFN1E1 \scheme[3]  (.D(\scheme_11[3] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[3]_net_1 ));
    DFN1E1 \randint[21]  (.D(\randint_12[21] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[21]_net_1 ));
    XOR2 un3_div_counter_I_7 (.A(N_5), .B(\div_counter[2]_net_1 ), .Y(
        I_7_0));
    NOR2A awaitscheme_RNO_3 (.A(N_500), .B(awaitheartbeat_net_1), .Y(
        awaitscheme_6_0_0_a3_0_0));
    OR3A awaitscheme_RNO_0 (.A(memo26), .B(N_309), .C(
        awaitscheme_6_0_0_o2_0), .Y(N_340));
    XOR2 un1_tick_3_I_26 (.A(\tick[0]_net_1 ), .B(N_336), .Y(
        \DWACT_ADD_CI_0_partial_sum[0] ));
    NOR2B un3_div_counter_I_6 (.A(\div_counter[1]_net_1 ), .B(
        \div_counter[0]_net_1 ), .Y(N_5));
    DFN1E1 \randint[3]  (.D(\randint_12[3] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[3]_net_1 ));
    DFN1 \counter[4]  (.D(\counter_17[4] ), .CLK(ref_signal_c), .Q(
        \counter[4]_net_1 ));
    NOR3A \frame_begin_RNO_1[2]  (.A(N_514), .B(\choice[2]_net_1 ), .C(
        \choice[1]_net_1 ), .Y(N_415));
    AX1 \cnt_RNO[3]  (.A(un1_start_1_sqmuxa_5), .B(cnt_c2), .C(
        cnt_n3_0), .Y(cnt_n3));
    AO13 \cnt_RNIOUCEK[1]  (.A(cnt_c0), .B(\cnt[1]_net_1 ), .C(
        cnt_0_sqmuxa), .Y(cnt_c1));
    DFN1E0C0 \data_size[4]  (.D(\data_size[3]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[4]_net_1 ));
    AO1A calculating_RNI78AS (.A(N_277), .B(calculating_net_1), .C(i44)
        , .Y(un1_i44));
    MX2 \scheme_RNO[24]  (.A(\scheme[30]_net_1 ), .B(
        demodulator_0_cur_scheme[24]), .S(init_2_net_1), .Y(
        \scheme_11[24] ));
    DFN1E0C0 \data_size[0]  (.D(\data_size[15]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[0]_net_1 ));
    XA1C \cnt_RNO[0]  (.A(cnt_n0_0_tz), .B(cnt_0_sqmuxa), .C(
        un1_start_1_sqmuxa_5), .Y(cnt_n0));
    AO1 calculating_RNIHA4RD (.A(un1_i44), .B(N_482), .C(
        start_1_sqmuxa), .Y(ilde_0_0_0));
    AO1 counting_RNO_0 (.A(un1_start_1_sqmuxa_1_0_0_a3_0), .B(N_443), 
        .C(start_1_sqmuxa), .Y(un1_start_1_sqmuxa_1_0_0_0));
    DFN1E1 choosing (.D(counting_0_sqmuxa_1), .CLK(ref_signal_c), .E(
        un1_counting_0_sqmuxa), .Q(choosing_net_1));
    DFN1E1 \scheme[41]  (.D(\scheme_11[41] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[41]_net_1 ));
    XOR3 un1_frame_begin_ADD_10x10_slow_I5_S (.A(\un1_choice_2[5] ), 
        .B(\frame_begin[5]_net_1 ), .C(I4_un1_CO1), .Y(
        \un1_frame_begin[5] ));
    OR3A launch_RNIIJ6R (.A(reset_c), .B(init_1_net_1), .C(
        launch_net_1), .Y(N_296));
    DFN1E1C0 \data_sent[9]  (.D(data_sent_n9), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[9]_net_1 ));
    XOR2 \data_sent_RNIVHFE[15]  (.A(\data_sent[15]_net_1 ), .B(
        \data_size[15]_net_1 ), .Y(un1_data_sent_15));
    NOR2 \div_counter_RNIL8VM[2]  (.A(\div_counter[2]_net_1 ), .B(
        \div_counter[3]_net_1 ), .Y(div_counter11_1));
    DFN1E1 \randint[17]  (.D(\randint_12[17] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[17]_net_1 ));
    DFN1E0C0 \data_size[2]  (.D(\data_size[1]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(N_14), .Q(
        \data_size[2]_net_1 ));
    NOR2B \flag_RNI9GN07[0]  (.A(cnt_0_sqmuxa_0), .B(counting_0_sqmuxa)
        , .Y(cnt_0_sqmuxa));
    AO1 \counter_RNO[5]  (.A(I_34), .B(un1_tick_2_sqmuxa_14), .C(N_505)
        , .Y(\counter_17[5] ));
    DFN1E1 head (.D(N_66), .CLK(ref_signal_c), .E(N_432), .Q(
        mac_0_head));
    OR2 start_RNI10BVT1 (.A(\tick_14_0_0_o2_2[4] ), .B(
        \tick_14_0_0_o2_1[4] ), .Y(N_320));
    XOR2 \data_sent_RNO[13]  (.A(data_sent_c12), .B(
        \data_sent[13]_net_1 ), .Y(data_sent_n13));
    XOR2 un1_tick_3_I_34 (.A(\tick[5]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12_1[0] ), .Y(I_34_0));
    NOR3C \data_sent_RNILF5I1[8]  (.A(\data_sent[7]_net_1 ), .B(
        data_sent_c6), .C(\data_sent[8]_net_1 ), .Y(data_sent_c8));
    NOR2A \data_len_RNO[3]  (.A(\scheme[0]_net_1 ), .B(
        demodulator_0_ctg[0]), .Y(\data_len_11[3] ));
    DFN1 \counter[1]  (.D(\counter_17[1] ), .CLK(ref_signal_c), .Q(
        \counter[1]_net_1 ));
    NOR3 \rd_RNI7F1F1[2]  (.A(\rd[0]_net_1 ), .B(\rd[2]_net_1 ), .C(
        \rd[1]_net_1 ), .Y(rd_0_sqmuxa_1_1));
    NOR2B \counter_RNO[0]  (.A(\DWACT_ADD_CI_0_partial_sum_0[0] ), .B(
        un1_tick_2_sqmuxa_14), .Y(\counter_17[0] ));
    OR2 resuming_RNO (.A(resuming_0_sqmuxa_2), .B(N_259), .Y(
        un1_resuming_0_sqmuxa_3));
    XO1 \data_size_RNICHUS[10]  (.A(\data_sent[10]_net_1 ), .B(
        \data_size[10]_net_1 ), .C(un1_data_sent_11), .Y(
        un1_data_sent_NE_1));
    MX2 \scheme_RNO[1]  (.A(\scheme[7]_net_1 ), .B(
        demodulator_0_cur_scheme[1]), .S(init_0_net_1), .Y(
        \scheme_11[1] ));
    XOR2 \data_size_RNIRDFE[13]  (.A(\data_size[13]_net_1 ), .B(
        \data_sent[13]_net_1 ), .Y(un1_data_sent_13));
    XAI1A \frame_begin_RNIQMJ7[9]  (.A(\counter[9]_net_1 ), .B(
        \frame_begin[9]_net_1 ), .C(awaitscheme7_2), .Y(blank17_NE_0));
    AND2 un1_tick_3_I_61 (.A(\DWACT_ADD_CI_0_pog_array_1_1[0] ), .B(
        \DWACT_ADD_CI_0_pog_array_1_2_0[0] ), .Y(
        \DWACT_ADD_CI_0_pog_array_2[0] ));
    XOR2 un1_counter_1_I_33 (.A(\counter[3]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12_0[0] ), .Y(I_33));
    MX2A \tick_RNO[2]  (.A(un1_tick_2_sqmuxa_2), .B(I_42_0), .S(N_213), 
        .Y(\tick_14[2] ));
    NOR2A calculating_RNIEBQRC (.A(N_283), .B(N_371), .Y(N_200));
    DFN1 \frame_begin[5]  (.D(N_48), .CLK(ref_signal_c), .Q(
        \frame_begin[5]_net_1 ));
    DFN1E1 \scheme[6]  (.D(\scheme_11[6] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[6]_net_1 ));
    XA1B \i_RNO[1]  (.A(\i[0]_net_1 ), .B(\i[1]_net_1 ), .C(
        un1_start_1_sqmuxa_7), .Y(N_874));
    NOR3 \counter_RNIF3682[5]  (.A(awaitscheme_6_0_0_o2_4_0), .B(
        awaitscheme_6_0_0_o2_4_1), .C(N_354), .Y(N_480));
    OA1 init_0_RNI7DURC2 (.A(N_464), .B(un1_tick_2_sqmuxa_10_1), .C(
        N_314), .Y(init_0_RNI7DURC2_net_1));
    AO1 sending_RNO_1 (.A(sending_7_i_i_a3_0_0), .B(N_276), .C(N_407), 
        .Y(sending_7_i_i_0));
    DFN1E1C0 \data_sent[6]  (.D(data_sent_n6), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[6]_net_1 ));
    NOR3A calculating_RNI9JOO6 (.A(un1_i44), .B(N_265), .C(N_269), .Y(
        i_1_sqmuxa));
    MX2 \scheme_RNO[5]  (.A(\scheme[11]_net_1 ), .B(
        demodulator_0_cur_scheme[5]), .S(init_0_net_1), .Y(
        \scheme_11[5] ));
    MX2 \scheme_RNO[3]  (.A(\scheme[9]_net_1 ), .B(
        demodulator_0_cur_scheme[3]), .S(init_0_net_1), .Y(
        \scheme_11[3] ));
    DFN1E1 \scheme[46]  (.D(N_348), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[46]_net_1 ));
    NOR2A \flag_RNIDUJD[0]  (.A(i44), .B(\flag[0]_net_1 ), .Y(N_487));
    NOR2B \rd_RNI35288[2]  (.A(rd_0_sqmuxa_1_1), .B(rd_0_sqmuxa), .Y(
        rd_0_sqmuxa_1));
    NOR3C \data_sent_RNIURMG[2]  (.A(\data_sent[0]_net_1 ), .B(
        \data_sent[1]_net_1 ), .C(\data_sent[2]_net_1 ), .Y(
        data_sent_c2));
    MAJ3 un1_frame_begin_ADD_10x10_slow_I4_un1_CO1 (.A(
        \frame_begin[4]_net_1 ), .B(N143), .C(\un1_choice_2[4] ), .Y(
        I4_un1_CO1));
    DFN1C0 \data_sent[0]  (.D(data_sent_e0), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\data_sent[0]_net_1 ));
    MX2 \randint_RNO[23]  (.A(\randint[2]_net_1 ), .B(
        randgen_0_cur_rand[23]), .S(init_1_net_1), .Y(\randint_12[23] )
        );
    DFN1E1 \data_len[7]  (.D(\data_len_11[7] ), .CLK(ref_signal_c), .E(
        un1_frame_begin_0_sqmuxa), .Q(\data_len[7]_net_1 ));
    MX2 \scheme_RNO[35]  (.A(\scheme[41]_net_1 ), .B(
        demodulator_0_cur_scheme[35]), .S(init_2_net_1), .Y(
        \scheme_11[35] ));
    MX2 \scheme_RNO[7]  (.A(\scheme[13]_net_1 ), .B(
        demodulator_0_cur_scheme[7]), .S(init_0_net_1), .Y(
        \scheme_11[7] ));
    OA1B \tick_RNIASN21[0]  (.A(\tick[1]_net_1 ), .B(\tick[0]_net_1 ), 
        .C(N_245), .Y(id_1_sqmuxa_1_i_0_a2_0));
    NOR2A \rd_RNO[2]  (.A(N_497), .B(rd_0_sqmuxa_1), .Y(\rd_13[2] ));
    MX2 \randint_RNO[17]  (.A(\randint[20]_net_1 ), .B(
        randgen_0_cur_rand[17]), .S(init_0_net_1), .Y(\randint_12[17] )
        );
    AX1 \cnt_RNO[2]  (.A(un1_start_1_sqmuxa_5), .B(cnt_c1), .C(
        cnt_n2_0), .Y(cnt_n2));
    DFN1E1 \randint[10]  (.D(\randint_12[10] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[10]_net_1 ));
    NOR3A counting_RNI4OL67 (.A(N_479), .B(N_281), .C(N_269), .Y(N_508)
        );
    NOR2B \choice_RNI6LOF7[1]  (.A(N_508), .B(\choice[1]_net_1 ), .Y(
        N_393));
    OR3 init_0_RNI0CAR91 (.A(N_505), .B(N_506), .C(un1_tick_2_sqmuxa_5)
        , .Y(un1_tick_2_sqmuxa_10_1));
    NOR2A \div_counter_RNO[5]  (.A(I_14_1), .B(div_counter11), .Y(
        \div_counter_3[5] ));
    DFN1 \counter[9]  (.D(\counter_17[9] ), .CLK(ref_signal_c), .Q(
        \counter[9]_net_1 ));
    NOR2B \tick_RNO[9]  (.A(I_38_0), .B(N_213), .Y(\tick_14[9] ));
    OR2 \tick_RNIG2Q6[9]  (.A(\tick[9]_net_1 ), .B(\tick[5]_net_1 ), 
        .Y(data_size_1_sqmuxa_i_0_o2_4_0));
    MX2 \scheme_RNO[41]  (.A(\scheme[47]_net_1 ), .B(
        demodulator_0_cur_scheme[41]), .S(init_net_1), .Y(
        \scheme_11[41] ));
    DFN1E1 \scheme[31]  (.D(\scheme_11[31] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[31]_net_1 ));
    NOR2B awaitbeacon_RNIJUM11 (.A(awaitbeacon_net_1), .B(N_245), .Y(
        N_456));
    XOR2 \memo_RNIEU6N[0]  (.A(\memo[0]_net_1 ), .B(
        demodulator_0_ord[0]), .Y(un1_ord_0));
    AX1C \data_sent_RNO[2]  (.A(\data_sent[0]_net_1 ), .B(
        \data_sent[1]_net_1 ), .C(\data_sent[2]_net_1 ), .Y(
        data_sent_n2));
    DFN1E1 launch (.D(un1_start_1_sqmuxa_6), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_4), .Q(launch_net_1));
    XO1 \data_size_RNIS1VS[14]  (.A(\data_sent[14]_net_1 ), .B(
        \data_size[14]_net_1 ), .C(un1_data_sent_15), .Y(
        un1_data_sent_NE_3));
    NOR2B \counter_RNO[8]  (.A(I_40), .B(un1_tick_2_sqmuxa_14), .Y(
        \counter_17[8] ));
    MX2 \scheme_RNO[17]  (.A(\scheme[23]_net_1 ), .B(
        demodulator_0_cur_scheme[17]), .S(init_2_net_1), .Y(
        \scheme_11[17] ));
    AND2 un1_tick_3_I_58 (.A(\tick[6]_net_1 ), .B(\tick[7]_net_1 ), .Y(
        \DWACT_ADD_CI_0_pog_array_1_2_0[0] ));
    XOR2 un1_rd_1_I_9 (.A(\rd[0]_net_1 ), .B(rd_0_sqmuxa), .Y(
        \DWACT_ADD_CI_0_partial_sum_1[0] ));
    NOR2A \tick_RNIQIGP[4]  (.A(sending13), .B(\tick[4]_net_1 ), .Y(
        un1_start_0_sqmuxa_0_0_a2_0_0));
    MAJ3 un1_frame_begin_ADD_10x10_slow_I6_un1_CO1 (.A(
        \frame_begin[6]_net_1 ), .B(N147), .C(\un1_choice_2[6] ), .Y(
        I6_un1_CO1));
    OA1C start_RNI78M5N (.A(start_net_1), .B(N_296), .C(
        un1_tick_2_sqmuxa_2), .Y(\tick_14_0_0_o2_2[4] ));
    DFN1 \tick[6]  (.D(\tick_14[6] ), .CLK(ref_signal_c), .Q(
        \tick[6]_net_1 ));
    NOR2B \tick_RNO[5]  (.A(I_34_0), .B(N_213), .Y(\tick_14[5] ));
    NOR2B \scheme_RNIV7HS7[2]  (.A(\scheme[2]_net_1 ), .B(N_474), .Y(
        \un1_choice_2[5] ));
    DFN1 \tick[1]  (.D(\tick_14[1] ), .CLK(ref_signal_c), .Q(
        \tick[1]_net_1 ));
    NOR3A calculating_RNISL0P6 (.A(rd_0_sqmuxa_0), .B(N_265), .C(N_269)
        , .Y(rd_0_sqmuxa));
    NOR3B start_RNIS6G46 (.A(N_476), .B(N_263), .C(N_276), .Y(
        un1_start_0_sqmuxa_0_0_a3_1));
    DFN1C0 \div_counter[1]  (.D(\div_counter_3[1] ), .CLK(ref_signal_c)
        , .CLR(reset_c), .Q(\div_counter[1]_net_1 ));
    NOR2 \choice_RNIFJ3O7[0]  (.A(\choice[0]_net_1 ), .B(N_284), .Y(
        N_514));
    DFN1E1 \scheme[5]  (.D(\scheme_11[5] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[5]_net_1 ));
    AO1 \tick_RNO_4[4]  (.A(N_478), .B(N_314), .C(I_35_0), .Y(N_358));
    NOR3A start_RNIHHDNB (.A(un1_tick_1_sqmuxa_2_i_i_a3_1), .B(N_299), 
        .C(sending_7_i_i_o2_0_1), .Y(N_432));
    OR2A init_1_RNIIVTAR (.A(N_338), .B(un1_tick_2_sqmuxa_5_0_0), .Y(
        un1_tick_2_sqmuxa_5));
    AO1A counting_RNIN4OUL (.A(N_259), .B(i_0_sqmuxa), .C(
        un1_start_1_sqmuxa_7_0_1_0), .Y(un1_start_1_sqmuxa_7));
    NOR2 \counter_RNIRO01[9]  (.A(\counter[9]_net_1 ), .B(
        \counter[6]_net_1 ), .Y(un1_tick_0_sqmuxa_1_0_a2_4_0));
    NOR2A \data_len_RNO[8]  (.A(\scheme[5]_net_1 ), .B(
        demodulator_0_ctg[0]), .Y(\data_len_11[8] ));
    AND2 un1_tick_3_I_59 (.A(\tick[2]_net_1 ), .B(\tick[3]_net_1 ), .Y(
        \DWACT_ADD_CI_0_pog_array_1[0] ));
    OR2 init_RNIQN6G4 (.A(N_329), .B(N_249), .Y(N_355));
    DFN1 \tick[7]  (.D(\tick_14[7] ), .CLK(ref_signal_c), .Q(
        \tick[7]_net_1 ));
    AX1C \data_sent_RNO[12]  (.A(\data_sent[11]_net_1 ), .B(
        data_sent_c10), .C(\data_sent[12]_net_1 ), .Y(data_sent_n12));
    AND2 un1_tick_3_I_1 (.A(\tick[0]_net_1 ), .B(N_336), .Y(
        \DWACT_ADD_CI_0_TMP[0] ));
    NOR3A choosing_RNINC8F1 (.A(N_472), .B(counting_net_1), .C(
        choosing_net_1), .Y(un1_calculating_0_sqmuxa_0_0_a3_0));
    DFN1E1 \scheme[43]  (.D(N_345), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[43]_net_1 ));
    DFN1E1 \scheme[36]  (.D(\scheme_11[36] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[36]_net_1 ));
    DFN1 \tick[0]  (.D(\tick_14[0] ), .CLK(ref_signal_c), .Q(
        \tick[0]_net_1 ));
    MX2 \flag_RNO[5]  (.A(\flag[6]_net_1 ), .B(
        demodulator_0_cur_flag[5]), .S(init_1_net_1), .Y(\flag_14[5] ));
    MX2 \scheme_RNO[21]  (.A(\scheme[27]_net_1 ), .B(
        demodulator_0_cur_scheme[21]), .S(init_2_net_1), .Y(
        \scheme_11[21] ));
    DFN1 \counter[5]  (.D(\counter_17[5] ), .CLK(ref_signal_c), .Q(
        \counter[5]_net_1 ));
    XO1 \data_size_RNIKPUS[12]  (.A(\data_sent[12]_net_1 ), .B(
        \data_size[12]_net_1 ), .C(un1_data_sent_13), .Y(
        un1_data_sent_NE_2));
    OR2A \i_RNI33FE[3]  (.A(\i[3]_net_1 ), .B(\i[2]_net_1 ), .Y(
        un1_resuming_0_sqmuxa_3_0_0_o3_0));
    DFN1E1 \scheme[15]  (.D(\scheme_11[15] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[15]_net_1 ));
    XOR2 un1_counter_1_I_40 (.A(\counter[8]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_3_0[0] ), .Y(I_40));
    MX2 \randint_RNO[18]  (.A(\randint[21]_net_1 ), .B(
        randgen_0_cur_rand[18]), .S(init_0_net_1), .Y(\randint_12[18] )
        );
    NOR3 calculating_RNI9JOO6_0 (.A(N_265), .B(N_269), .C(un1_i44), .Y(
        i_0_sqmuxa));
    OA1 init_1_RNI361P6 (.A(N_274), .B(N_249), .C(init_1_net_1), .Y(
        N_42));
    XA1C \cnt_RNO_1[3]  (.A(\cnt[3]_net_1 ), .B(cnt_0_sqmuxa), .C(
        un1_start_1_sqmuxa_5), .Y(cnt_n3_0));
    AND2 un1_counter_1_I_1 (.A(\counter[0]_net_1 ), .B(
        init_0_RNI7DURC2_net_1), .Y(\DWACT_ADD_CI_0_TMP_0[0] ));
    DFN1E1 \scheme[17]  (.D(\scheme_11[17] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[17]_net_1 ));
    NOR2A \tick_RNIM924D[4]  (.A(data_sent_1_sqmuxa_1_1), .B(N_355), 
        .Y(data_sent_1_sqmuxa_1));
    NOR2B \counter_RNO[4]  (.A(I_35), .B(un1_tick_2_sqmuxa_14), .Y(
        \counter_17[4] ));
    DFN1E1 \scheme[25]  (.D(\scheme_11[25] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[25]_net_1 ));
    DFN1E1 \data_len[8]  (.D(\data_len_11[8] ), .CLK(ref_signal_c), .E(
        un1_frame_begin_0_sqmuxa), .Q(\data_len[8]_net_1 ));
    OR2A launch_RNO_0 (.A(N_200), .B(un1_start_1_sqmuxa_4_0), .Y(
        un1_start_1_sqmuxa_4));
    NOR2B \tick_RNO[7]  (.A(I_39_0), .B(N_213), .Y(\tick_14[7] ));
    OR3A \tick_RNI6H6A[2]  (.A(\tick[2]_net_1 ), .B(\tick[1]_net_1 ), 
        .C(\tick[0]_net_1 ), .Y(N_278));
    DFN1E1 \scheme[40]  (.D(\scheme_11[40] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[40]_net_1 ));
    AX1C \data_sent_RNO[8]  (.A(\data_sent[7]_net_1 ), .B(data_sent_c6)
        , .C(\data_sent[8]_net_1 ), .Y(data_sent_n8));
    XOR2 \cnt_RNO_0[1]  (.A(cnt_c0), .B(\cnt[1]_net_1 ), .Y(
        cnt_n1_0_tz));
    MX2 \scheme_RNO[10]  (.A(\scheme[16]_net_1 ), .B(
        demodulator_0_cur_scheme[10]), .S(init_1_net_1), .Y(
        \scheme_11[10] ));
    NOR2B calculating_RNIBLML7 (.A(i_0_sqmuxa), .B(N_259), .Y(
        flag_1_sqmuxa));
    DFN1E1 \scheme[27]  (.D(\scheme_11[27] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[27]_net_1 ));
    NOR2A \rd_RNO[0]  (.A(N_495), .B(rd_0_sqmuxa_1), .Y(\rd_13[0] ));
    XOR2 un1_tick_3_I_40 (.A(\tick[8]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_3[0] ), .Y(I_40_0));
    OR3 \tick_RNIC3EK[3]  (.A(data_size_1_sqmuxa_i_0_o2_4_1), .B(
        data_size_1_sqmuxa_i_0_o2_4_0), .C(
        data_size_1_sqmuxa_i_0_o2_4_2), .Y(N_268));
    OR3 \data_size_RNI4VD33[12]  (.A(un1_data_sent_NE_3), .B(
        un1_data_sent_NE_2), .C(un1_data_sent_NE_8), .Y(
        un1_data_sent_NE_12));
    NOR2A blank_RNILIHB9 (.A(start_2_sqmuxa), .B(blank18), .Y(
        start_0_sqmuxa));
    XO1 \data_size_RNI0AHC[6]  (.A(\data_sent[6]_net_1 ), .B(
        \data_size[6]_net_1 ), .C(un1_data_sent_7), .Y(
        un1_data_sent_NE_7));
    NOR2A \data_len_RNO[4]  (.A(\scheme[1]_net_1 ), .B(
        demodulator_0_ctg[0]), .Y(\data_len_11[4] ));
    OR2A \tick_RNIBG9T1[4]  (.A(N_288), .B(N_478), .Y(
        data_size_1_sqmuxa_i_0_0));
    NOR2A \randint_RNO[11]  (.A(\randint[14]_net_1 ), .B(init_net_1), 
        .Y(\randint_12[11] ));
    NOR2 \i_RNO[0]  (.A(un1_start_1_sqmuxa_7), .B(\i[0]_net_1 ), .Y(
        N_873));
    XA1B \frame_begin_RNO[7]  (.A(I6_un1_CO1), .B(
        ADD_10x10_slow_I7_S_0), .C(N_63), .Y(\frame_begin_18[7] ));
    NOR3B \counter_RNI7DTF1[5]  (.A(un1_tick_0_sqmuxa_1_0_a2_4_0), .B(
        un1_tick_0_sqmuxa_1_0_a2_4_1), .C(N_265), .Y(N_477));
    NOR2B \cnt_RNI1NPF6[3]  (.A(resuming_0_sqmuxa_2_0_a2_0_a3_2), .B(
        resuming_0_sqmuxa), .Y(resuming_0_sqmuxa_2));
    MX2 \scheme_RNO[29]  (.A(\scheme[35]_net_1 ), .B(
        demodulator_0_cur_scheme[29]), .S(init_2_net_1), .Y(
        \scheme_11[29] ));
    NOR2A resuming_RNIDF1C (.A(resuming_net_1), .B(counting_net_1), .Y(
        tick_1_sqmuxa_3_i_i_a3_0));
    NOR3B init_0_RNIC1VK3 (.A(un1_tick_2_sqmuxa_5_0_a2_1), .B(
        div_counter11), .C(init_0_net_1), .Y(
        un1_tick_2_sqmuxa_5_0_a2_3));
    XOR2 \data_size_RNITH86[5]  (.A(\data_size[5]_net_1 ), .B(
        \data_sent[5]_net_1 ), .Y(un1_data_sent_5));
    NOR2B \tick_RNO[0]  (.A(\DWACT_ADD_CI_0_partial_sum[0] ), .B(N_213)
        , .Y(\tick_14[0] ));
    DFN1E1C0 sending (.D(N_158), .CLK(ref_signal_c), .CLR(reset_c), .E(
        div_counter11), .Q(mac_0_sending));
    NOR2A choosing_RNITTL6 (.A(choosing_net_1), .B(counting_net_1), .Y(
        i44));
    NOR2B \choice_RNI7MOF7[2]  (.A(N_508), .B(\choice[2]_net_1 ), .Y(
        N_434));
    OR2A \counter_RNINK01[5]  (.A(\counter[6]_net_1 ), .B(
        \counter[5]_net_1 ), .Y(awaitscheme_6_0_0_o2_4_1));
    OR2 blank_RNIVE7F (.A(blank_net_1), .B(launch_net_1), .Y(N_264));
    NOR2A \randint_RNO[0]  (.A(\randint[3]_net_1 ), .B(init_net_1), .Y(
        \randint_12[0] ));
    NOR3C \data_sent_RNIKF071[6]  (.A(\data_sent[5]_net_1 ), .B(
        data_sent_c4), .C(\data_sent[6]_net_1 ), .Y(data_sent_c6));
    OR2 awaitscheme_RNIKURD1 (.A(N_252), .B(N_245), .Y(N_265));
    NOR2B un1_frame_begin_ADD_10x10_slow_I2_un3_CO1 (.A(N_378), .B(
        \frame_begin[2]_net_1 ), .Y(I2_un1_CO1));
    MX2 \scheme_RNO[28]  (.A(\scheme[34]_net_1 ), .B(
        demodulator_0_cur_scheme[28]), .S(init_2_net_1), .Y(
        \scheme_11[28] ));
    NOR2B un1_tick_3_I_53 (.A(\DWACT_ADD_CI_0_g_array_2[0] ), .B(
        \DWACT_ADD_CI_0_pog_array_2[0] ), .Y(
        \DWACT_ADD_CI_0_g_array_3[0] ));
    DFN1E1 \scheme[33]  (.D(\scheme_11[33] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[33]_net_1 ));
    MX2 \randint_RNO[22]  (.A(\randint[1]_net_1 ), .B(
        randgen_0_cur_rand[22]), .S(init_1_net_1), .Y(\randint_12[22] )
        );
    NOR3B \counter_RNIQLVT[5]  (.A(un1_tick_0_sqmuxa_1_0_a2_4_0), .B(
        un1_tick_0_sqmuxa_1_0_a2_4_1), .C(N_245), .Y(N_500));
    DFN1C0 awaitheartbeat (.D(awaitheartbeat_RNO_net_1), .CLK(
        ref_signal_c), .CLR(reset_c), .Q(awaitheartbeat_net_1));
    NOR2A \data_len_RNO[5]  (.A(\scheme[2]_net_1 ), .B(
        demodulator_0_ctg[0]), .Y(\data_len_11[5] ));
    AO1 \counter_RNO[6]  (.A(I_36), .B(un1_tick_2_sqmuxa_14), .C(N_506)
        , .Y(\counter_17[6] ));
    XOR2 un1_tick_3_I_38 (.A(\tick[9]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12_3[0] ), .Y(I_38_0));
    NOR2A resuming_RNIQEI81 (.A(resuming_net_1), .B(N_259), .Y(N_472));
    NOR2B \tick_RNO[8]  (.A(I_40_0), .B(N_213), .Y(\tick_14[8] ));
    NOR3C resuming_RNIUS327 (.A(N_259), .B(resuming_net_1), .C(N_481), 
        .Y(N_400));
    NOR2B \scheme_RNI1AHS7[4]  (.A(\scheme[4]_net_1 ), .B(N_474), .Y(
        \un1_choice_2[7] ));
    NOR3B start_RNIDCQ53 (.A(div_counter11), .B(start_net_1), .C(N_296)
        , .Y(un1_tick_1_sqmuxa_2_i_i_a3_1));
    MX2 \scheme_RNO[12]  (.A(\scheme[18]_net_1 ), .B(
        demodulator_0_cur_scheme[12]), .S(init_1_net_1), .Y(
        \scheme_11[12] ));
    NOR3B head_RNO_2 (.A(N_245), .B(N_325), .C(\id[2]_net_1 ), .Y(
        N_384));
    AO1 \counter_RNO[9]  (.A(I_38), .B(un1_tick_2_sqmuxa_14), .C(N_506)
        , .Y(\counter_17[9] ));
    OR2 awaitbeacon_RNI0J5J (.A(awaitbeacon_net_1), .B(
        awaitheartbeat_net_1), .Y(awaitscheme_6_0_0_o2_0_0));
    MX2 \scheme_RNO[13]  (.A(\scheme[19]_net_1 ), .B(
        demodulator_0_cur_scheme[13]), .S(init_1_net_1), .Y(
        \scheme_11[13] ));
    XOR2 un1_tick_3_I_39 (.A(\tick[7]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12_2[0] ), .Y(I_39_0));
    DFN1E1 \randint[6]  (.D(\randint_12[6] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[6]_net_1 ));
    DFN1E1C0 \data_sent[7]  (.D(data_sent_n7), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[7]_net_1 ));
    DFN1E1 \scheme[30]  (.D(\scheme_11[30] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[30]_net_1 ));
    DFN1E1 \randint[15]  (.D(\randint_12[15] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[15]_net_1 ));
    XO1 \frame_begin_RNI426D[4]  (.A(\frame_begin[4]_net_1 ), .B(
        \counter[4]_net_1 ), .C(blank17_3), .Y(blank17_NE_2));
    AND3 un3_div_counter_I_10 (.A(\div_counter[0]_net_1 ), .B(
        \div_counter[1]_net_1 ), .C(\div_counter[2]_net_1 ), .Y(
        \DWACT_FINC_E[0] ));
    DFN1E1C0 \memo[1]  (.D(demodulator_0_ord[1]), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(N_149), .Q(\memo[1]_net_1 ));
    DFN1E1 \randint[11]  (.D(\randint_12[11] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[11]_net_1 ));
    AX1C \data_sent_RNO[6]  (.A(\data_sent[5]_net_1 ), .B(data_sent_c4)
        , .C(\data_sent[6]_net_1 ), .Y(data_sent_n6));
    OR2 blank_RNO_0 (.A(start_0_sqmuxa), .B(start_1_sqmuxa), .Y(
        un1_tick_2_sqmuxa_0));
    NOR3A sending_RNO_4 (.A(start_net_1), .B(init_0_net_1), .C(
        launch_net_1), .Y(sending_7_i_i_a3_2_0));
    DFN1 \cnt[1]  (.D(cnt_n1), .CLK(ref_signal_c), .Q(\cnt[1]_net_1 ));
    OR2A launch_RNINJR7L (.A(N_200), .B(tick_2_sqmuxa), .Y(N_464));
    NOR3A choosing_RNILAAI_0 (.A(resuming_net_1), .B(counting_net_1), 
        .C(choosing_net_1), .Y(N_395_1));
    NOR2B un1_tick_3_I_47 (.A(\DWACT_ADD_CI_0_g_array_2[0] ), .B(
        \tick[4]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12_1[0] ));
    NOR2A \div_counter_RNIH4VM[1]  (.A(\div_counter[0]_net_1 ), .B(
        \div_counter[1]_net_1 ), .Y(div_counter11_2));
    XOR2 un1_rd_1_I_12 (.A(\DWACT_ADD_CI_0_partial_sum[1] ), .B(
        \DWACT_ADD_CI_0_TMP_1[0] ), .Y(I_12_0));
    XA1B \frame_begin_RNO[9]  (.A(\frame_begin[9]_net_1 ), .B(
        I8_un1_CO1), .C(N_63), .Y(\frame_begin_18[9] ));
    XOR2 \choice_RNI0BAG[0]  (.A(\choice[0]_net_1 ), .B(\i[0]_net_1 ), 
        .Y(N_248_i));
    DFN1E1 \randint[7]  (.D(\randint_12[7] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[7]_net_1 ));
    MX2 \scheme_RNO[16]  (.A(\scheme[22]_net_1 ), .B(
        demodulator_0_cur_scheme[16]), .S(init_1_net_1), .Y(
        \scheme_11[16] ));
    DFN1 \frame_begin[6]  (.D(N_46), .CLK(ref_signal_c), .Q(
        \frame_begin[6]_net_1 ));
    NOR2B init_0_RNIBHAK7 (.A(N_483), .B(N_480), .Y(N_506));
    NOR2 \data_len_RNI7SB7[5]  (.A(\data_len[5]_net_1 ), .B(
        \data_len[6]_net_1 ), .Y(sending13_2));
    MX2 \randint_RNO[14]  (.A(\randint[17]_net_1 ), .B(
        randgen_0_cur_rand[14]), .S(init_0_net_1), .Y(\randint_12[14] )
        );
    NOR3 working_RNO (.A(N_411), .B(N_410), .C(N_409), .Y(N_55));
    NOR2A \randint_RNO[4]  (.A(\randint[7]_net_1 ), .B(init_net_1), .Y(
        \randint_12[4] ));
    XA1C \cnt_RNO_0[2]  (.A(\cnt[2]_net_1 ), .B(cnt_0_sqmuxa), .C(
        un1_start_1_sqmuxa_5), .Y(cnt_n2_0));
    XOR2 un1_tick_3_I_42 (.A(\tick[2]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_1[0] ), .Y(I_42_0));
    DFN1E1 \scheme[19]  (.D(\scheme_11[19] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[19]_net_1 ));
    XOR2 un1_frame_begin_ADD_10x10_slow_I3_S_0 (.A(
        \frame_begin[3]_net_1 ), .B(I2_un1_CO1), .Y(
        ADD_10x10_slow_I3_S_0));
    MX2 \randint_RNO[13]  (.A(\randint[16]_net_1 ), .B(
        randgen_0_cur_rand[13]), .S(init_0_net_1), .Y(\randint_12[13] )
        );
    NOR2A \data_len_RNO[7]  (.A(\scheme[4]_net_1 ), .B(
        demodulator_0_ctg[0]), .Y(\data_len_11[7] ));
    DFN1E1 calculating (.D(calculating_0_sqmuxa), .CLK(ref_signal_c), 
        .E(un1_calculating_0_sqmuxa), .Q(calculating_net_1));
    OR3 awaitbeacon_RNISK462 (.A(N_504), .B(awaitbeacon_net_1), .C(
        N_244), .Y(N_354));
    NOR2B un1_counter_1_I_44 (.A(\DWACT_ADD_CI_0_g_array_3_0[0] ), .B(
        \counter[8]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12_3_0[0] ));
    DFN1 \tick[2]  (.D(\tick_14[2] ), .CLK(ref_signal_c), .Q(
        \tick[2]_net_1 ));
    OR2 \frame_begin_RNO_0[4]  (.A(N_505), .B(N_514), .Y(
        \frame_begin_18_i_0_0[4] ));
    NOR2B un1_counter_1_I_55 (.A(\DWACT_ADD_CI_0_g_array_1_0[0] ), .B(
        \DWACT_ADD_CI_0_pog_array_1_0[0] ), .Y(
        \DWACT_ADD_CI_0_g_array_2_0[0] ));
    OR3 \data_size_RNIGM3I1[0]  (.A(un1_data_sent_NE_5), .B(
        un1_data_sent_NE_4), .C(un1_data_sent_NE_11), .Y(
        un1_data_sent_NE_13));
    DFN1E1 \scheme[29]  (.D(\scheme_11[29] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[29]_net_1 ));
    OA1C \frame_begin_RNO[4]  (.A(N_284), .B(\un1_frame_begin[4] ), .C(
        \frame_begin_18_i_0_0[4] ), .Y(N_50));
    OA1 resuming_RNIHTI56 (.A(counting_net_1), .B(resuming_net_1), .C(
        N_481), .Y(N_423));
    DFN1E0C0 \id[0]  (.D(\id[2]_net_1 ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_16), .Q(\id[0]_net_1 ));
    NOR3A calculating_RNO (.A(un1_calculating_0_sqmuxa_0_0_a3_0), .B(
        N_265), .C(N_269), .Y(calculating_0_sqmuxa));
    XOR2 \data_sent_RNO[14]  (.A(data_sent_c13), .B(
        \data_sent[14]_net_1 ), .Y(data_sent_n14));
    AO1 init_0_RNIT1GFJ (.A(blank18), .B(start_2_sqmuxa), .C(N_154), 
        .Y(un1_tick_2_sqmuxa_5_0_0));
    AO1A \tick_RNIF4UG4[4]  (.A(N_354), .B(
        un1_start_0_sqmuxa_0_0_a2_0_0), .C(N_458), .Y(N_263));
    XOR2 un1_rd_1_I_7 (.A(\rd[1]_net_1 ), .B(rd_0_sqmuxa), .Y(
        \DWACT_ADD_CI_0_pog_array_0[0] ));
    MX2 \randint_RNO[16]  (.A(\randint[19]_net_1 ), .B(
        randgen_0_cur_rand[16]), .S(init_0_net_1), .Y(\randint_12[16] )
        );
    DFN1E1 \data_len[6]  (.D(\data_len_11[6] ), .CLK(ref_signal_c), .E(
        un1_frame_begin_0_sqmuxa), .Q(\data_len[6]_net_1 ));
    XOR2 un1_counter_1_I_26 (.A(\counter[0]_net_1 ), .B(
        init_0_RNI7DURC2_net_1), .Y(\DWACT_ADD_CI_0_partial_sum_0[0] ));
    DFN1C0 \div_counter[0]  (.D(I_4_0), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\div_counter[0]_net_1 ));
    OR2 \i_RNIVUEE_0[1]  (.A(\i[1]_net_1 ), .B(\i[0]_net_1 ), .Y(N_256)
        );
    DFN1 \cnt[2]  (.D(cnt_n2), .CLK(ref_signal_c), .Q(\cnt[2]_net_1 ));
    XO1 \frame_begin_RNICA6D[5]  (.A(\frame_begin[5]_net_1 ), .B(
        \counter[5]_net_1 ), .C(blank17_6), .Y(blank17_NE_3));
    DFN1E1 \flag[3]  (.D(\flag_14[3] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_2), .Q(\flag[3]_net_1 ));
    DFN1 \counter[8]  (.D(\counter_17[8] ), .CLK(ref_signal_c), .Q(
        \counter[8]_net_1 ));
    OR2 awaitscheme_RNIDNTH (.A(awaitscheme_net_1), .B(
        awaitheartbeat_net_1), .Y(N_252));
    NOR3A resuming_RNO_1 (.A(N_395_1), .B(N_265), .C(N_269), .Y(N_386));
    MX2 \scheme_RNO[14]  (.A(\scheme[20]_net_1 ), .B(
        demodulator_0_cur_scheme[14]), .S(init_1_net_1), .Y(
        \scheme_11[14] ));
    MX2 \randint_RNO[6]  (.A(\randint[9]_net_1 ), .B(
        randgen_0_cur_rand[6]), .S(init_net_1), .Y(\randint_12[6] ));
    XOR2 \data_sent_RNO[1]  (.A(\data_sent[1]_net_1 ), .B(
        \data_sent[0]_net_1 ), .Y(data_sent_n1));
    DFN1E1 \data_len[5]  (.D(\data_len_11[5] ), .CLK(ref_signal_c), .E(
        un1_frame_begin_0_sqmuxa), .Q(\data_len[5]_net_1 ));
    OA1C \frame_begin_RNO[6]  (.A(N_284), .B(\un1_frame_begin[6] ), .C(
        \frame_begin_18_i_0_0[6] ), .Y(N_46));
    DFN1E1 \randint[16]  (.D(\randint_12[16] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa), .Q(\randint[16]_net_1 ));
    OR3 choosing_RNILAAI (.A(counting_net_1), .B(resuming_net_1), .C(
        choosing_net_1), .Y(N_277));
    MX2 \scheme_RNO[45]  (.A(\scheme[3]_net_1 ), .B(
        demodulator_0_cur_scheme[45]), .S(init_net_1), .Y(N_347));
    VCC VCC_i (.Y(VCC));
    XOR2 un1_tick_3_I_33 (.A(\tick[3]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12[0] ), .Y(I_33_0));
    OR3 resuming_RNIBRFPQ (.A(ilde_0_0_0), .B(N_423), .C(i_0_sqmuxa), 
        .Y(ie));
    OR2 init_RNITUQS (.A(N_276), .B(init_net_1), .Y(N_329));
    XOR2 \frame_begin_RNI98J6[7]  (.A(\counter[7]_net_1 ), .B(
        \frame_begin[7]_net_1 ), .Y(blank17_7));
    NOR2B init_0_RNI3R1S6 (.A(N_483), .B(N_477), .Y(N_505));
    NOR2A \flag_RNII2S31[0]  (.A(N_259), .B(\flag[0]_net_1 ), .Y(
        cnt_0_sqmuxa_0));
    XO1 \choice_RNI4QK01[2]  (.A(\i[2]_net_1 ), .B(\choice[2]_net_1 ), 
        .C(N_248_i), .Y(un1_resuming_0_sqmuxa_5_0_0_o2_1));
    DFN1E1C0 awaitscheme (.D(awaitscheme_6), .CLK(ref_signal_c), .CLR(
        reset_c), .E(div_counter11), .Q(awaitscheme_net_1));
    XOR2 un1_frame_begin_ADD_10x10_slow_I8_S_0 (.A(
        \frame_begin[8]_net_1 ), .B(\un1_choice_2[8] ), .Y(
        ADD_10x10_slow_I8_S_0));
    OR3A blank_RNIQNKP61 (.A(N_314), .B(N_249), .C(N_461), .Y(
        \tick_14_0_0_o2_1[4] ));
    NOR2B un1_tick_3_I_56 (.A(\DWACT_ADD_CI_0_TMP[0] ), .B(
        \tick[1]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_1[0] ));
    XOR2 un1_counter_1_I_34 (.A(\counter[5]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12_1_0[0] ), .Y(I_34));
    XOR2 un1_counter_1_I_42 (.A(\counter[2]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_1_0[0] ), .Y(I_42));
    NOR3 \i_RNIFJA73[3]  (.A(un1_resuming_0_sqmuxa_5_0_0_o2_0), .B(
        un1_resuming_0_sqmuxa_5_0_0_o2_1), .C(N_281), .Y(
        un1_resuming_0_sqmuxa_5_0_0_a2_0));
    AO1D \frame_begin_RNO_0[5]  (.A(\choice[1]_net_1 ), .B(N_284), .C(
        N_505), .Y(\frame_begin_18_i_0_0[5] ));
    DFN1 \frame_begin[7]  (.D(\frame_begin_18[7] ), .CLK(ref_signal_c), 
        .Q(\frame_begin[7]_net_1 ));
    DFN1 \rd[0]  (.D(\rd_13[0] ), .CLK(ref_signal_c), .Q(\rd[0]_net_1 )
        );
    NOR2B \flag_RNIUGT56[0]  (.A(N_487), .B(N_482), .Y(N_396));
    NOR3C \data_sent_RNINJRR[4]  (.A(\data_sent[3]_net_1 ), .B(
        data_sent_c2), .C(\data_sent[4]_net_1 ), .Y(data_sent_c4));
    AND2 un1_counter_1_I_60 (.A(\counter[4]_net_1 ), .B(
        \counter[5]_net_1 ), .Y(\DWACT_ADD_CI_0_pog_array_1_1_0[0] ));
    DFN1E1 past (.D(un1_tick_0_sqmuxa), .CLK(ref_signal_c), .E(
        un1_tick_0_sqmuxa_1), .Q(past_net_1));
    DFN1E1 \scheme[12]  (.D(\scheme_11[12] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[12]_net_1 ));
    DFN1E0P0 \data_size[3]  (.D(\data_size[2]_net_1 ), .CLK(
        ref_signal_c), .PRE(reset_c), .E(N_14), .Q(
        \data_size[3]_net_1 ));
    OR2 start_RNO (.A(un1_tick_0_sqmuxa_1_1_0), .B(start_0_sqmuxa), .Y(
        un1_start_0_sqmuxa));
    DFN1 \tick[9]  (.D(\tick_14[9] ), .CLK(ref_signal_c), .Q(
        \tick[9]_net_1 ));
    NOR2A \rd_RNO[1]  (.A(N_496), .B(rd_0_sqmuxa_1), .Y(\rd_13[1] ));
    MAJ3 un1_frame_begin_ADD_10x10_slow_I8_un1_CO1 (.A(
        \frame_begin[8]_net_1 ), .B(N151), .C(\un1_choice_2[8] ), .Y(
        I8_un1_CO1));
    DFN1E1 \scheme[22]  (.D(\scheme_11[22] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[22]_net_1 ));
    XOR2 un1_counter_1_I_39 (.A(\counter[7]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12_2_0[0] ), .Y(I_39));
    OR3 \frame_begin_RNITJPL1[4]  (.A(blank17_NE_2), .B(blank17_NE_1), 
        .C(blank17_NE_6), .Y(blank18));
    NOR2B \tick_RNO[1]  (.A(I_37_0), .B(N_213), .Y(\tick_14[1] ));
    NOR2 \i_RNIGDOOD_0[1]  (.A(N_200), .B(N_259), .Y(N_444));
    OA1C \tick_RNO_5[4]  (.A(N_252), .B(N_449), .C(awaitbeacon_net_1), 
        .Y(\tick_14_0_0_a3_2_2_0[4] ));
    XOR2 \frame_begin_RNIVTI6[2]  (.A(\counter[2]_net_1 ), .B(
        \frame_begin[2]_net_1 ), .Y(blank17_2));
    DFN1E1 \scheme[45]  (.D(N_347), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[45]_net_1 ));
    DFN1E1 \scheme[1]  (.D(\scheme_11[1] ), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3_0), .Q(\scheme[1]_net_1 ));
    DFN1C0 \div_counter[2]  (.D(I_7_0), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\div_counter[2]_net_1 ));
    DFN1E1C0 \data_sent[1]  (.D(data_sent_n1), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(data_sent_1_sqmuxa_1), .Q(
        \data_sent[1]_net_1 ));
    DFN1E0P0 \data_size[1]  (.D(\data_size[0]_net_1 ), .CLK(
        ref_signal_c), .PRE(reset_c), .E(N_14), .Q(
        \data_size[1]_net_1 ));
    MX2 \scheme_RNO[25]  (.A(\scheme[31]_net_1 ), .B(
        demodulator_0_cur_scheme[25]), .S(init_2_net_1), .Y(
        \scheme_11[25] ));
    AO1D head_RNO_0 (.A(N_361), .B(N_245), .C(N_384), .Y(head_13_0_i_0)
        );
    XOR2 un3_div_counter_I_9 (.A(N_4), .B(\div_counter[3]_net_1 ), .Y(
        I_9_0));
    MX2 \flag_RNO[7]  (.A(\flag[0]_net_1 ), .B(
        demodulator_0_cur_flag[7]), .S(init_1_net_1), .Y(\flag_14[7] ));
    DFN1E1 \scheme[47]  (.D(N_349), .CLK(ref_signal_c), .E(
        un1_start_1_sqmuxa_3), .Q(\scheme[47]_net_1 ));
    
endmodule


module modulator(
       reset_c,
       ref_signal_c,
       trigger_signal_c,
       output_signal_c
    );
input  reset_c;
input  ref_signal_c;
input  trigger_signal_c;
output output_signal_c;

    wire output_signal_0, output_signal_1_sqmuxa_i_3, 
        output_signal_1_sqmuxa_i_1, N_147, N_148, 
        \clock_counter[14]_net_1 , \clock_counter[15]_net_1 , N_36_3, 
        output_signal_1_sqmuxa_i_a2_2, output_signal_1_sqmuxa_i_a2_1, 
        \clock_counter[9]_net_1 , \clock_counter[10]_net_1 , un6lto11, 
        un6lto12, output_signal_1_sqmuxa_i_a2_0_2, 
        \clock_counter[8]_net_1 , \clock_counter[6]_net_1 , 
        output_signal_1_sqmuxa_i_a2_0_1, \clock_counter[5]_net_1 , 
        \clock_counter[4]_net_1 , counter_n1_i_0, \counter[0]_net_1 , 
        \counter[1]_net_1 , output_signal_1_sqmuxa_i_a2_3_0, 
        output_signal_1_sqmuxa_i_a2_2_0, un6lto7, 
        counter_0_sqmuxa_i_a2_0, N_123_1, clock_counterlde_0_a2_1, 
        \counter[4]_net_1 , \counter[5]_net_1 , 
        output_signal_1_sqmuxa_i_o2_0, \clock_counter[2]_net_1 , 
        \clock_counter[3]_net_1 , N_5, N_151, \counter[2]_net_1 , 
        \counter[3]_net_1 , N_19, N_53, counter_n0, N_21, N_139, N_23, 
        N_42, N_25, N_41, N_27, N_40, N_29, N_39, N_31, 
        \clock_counter[0]_net_1 , \clock_counter[1]_net_1 , N_17, N_46, 
        N_137, N_150, N_55, N_145, N_45, N_146, N_47, N_36, N_51, 
        counter_n2, counter_c1, N_8, counter_n3, counter_c2, 
        counter_n5, counter_44_0, counter_n4, counter_c3, N_144, 
        clock_countere, \clock_counter[13]_net_1 , N_91, N_52, N_61, 
        N_50, N_49, N_48, clock_counter_n9, clock_counter_n10, 
        clock_counter_n11, clock_counter_n12, clock_counter_n13, 
        clock_counter_n14, clock_counter_n15, GND, VCC;
    
    OR2 \clock_counter_RNIJ3G2[2]  (.A(\clock_counter[2]_net_1 ), .B(
        \clock_counter[3]_net_1 ), .Y(output_signal_1_sqmuxa_i_o2_0));
    DFN1E1C0 \clock_counter[6]  (.D(N_21), .CLK(ref_signal_c), .CLR(
        reset_c), .E(clock_countere), .Q(\clock_counter[6]_net_1 ));
    XA1A \clock_counter_RNO[4]  (.A(\clock_counter[4]_net_1 ), .B(N_41)
        , .C(counter_n0), .Y(N_25));
    NOR2B \counter_RNINTKF1[2]  (.A(counter_c1), .B(\counter[2]_net_1 )
        , .Y(counter_c2));
    DFN1E1C0 \clock_counter[3]  (.D(N_27), .CLK(ref_signal_c), .CLR(
        reset_c), .E(clock_countere), .Q(\clock_counter[3]_net_1 ));
    NOR3 \counter_RNIT3LF1[5]  (.A(\counter[4]_net_1 ), .B(
        \counter[5]_net_1 ), .C(\counter[0]_net_1 ), .Y(
        clock_counterlde_0_a2_1));
    DFN1E1C0 \clock_counter[4]  (.D(N_25), .CLK(ref_signal_c), .CLR(
        reset_c), .E(clock_countere), .Q(\clock_counter[4]_net_1 ));
    DFN1E1C0 \clock_counter[8]  (.D(N_17), .CLK(ref_signal_c), .CLR(
        reset_c), .E(clock_countere), .Q(\clock_counter[8]_net_1 ));
    DFN1C0 \counter[2]  (.D(counter_n2), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[2]_net_1 ));
    DFN1E1C0 \clock_counter[1]  (.D(N_31), .CLK(ref_signal_c), .CLR(
        reset_c), .E(clock_countere), .Q(\clock_counter[1]_net_1 ));
    DFN1E1C0 \clock_counter[0]  (.D(N_144), .CLK(ref_signal_c), .CLR(
        reset_c), .E(clock_countere), .Q(\clock_counter[0]_net_1 ));
    NOR2A output_signal_RNO_7 (.A(output_signal_1_sqmuxa_i_a2_3_0), .B(
        N_55), .Y(N_150));
    OR3B \clock_counter_RNI6GO8[6]  (.A(\clock_counter[5]_net_1 ), .B(
        \clock_counter[6]_net_1 ), .C(N_42), .Y(N_53));
    OR2A \clock_counter_RNI2305[3]  (.A(\clock_counter[3]_net_1 ), .B(
        N_40), .Y(N_41));
    OR2A \clock_counter_RNI41VU[11]  (.A(un6lto11), .B(N_48), .Y(N_49));
    XA1B \counter_RNO[4]  (.A(\counter[4]_net_1 ), .B(counter_c3), .C(
        N_8), .Y(counter_n4));
    OR2A \clock_counter_RNID686[4]  (.A(\clock_counter[4]_net_1 ), .B(
        N_41), .Y(N_42));
    VCC VCC_i (.Y(VCC));
    NOR2A \clock_counter_RNO[0]  (.A(counter_n0), .B(
        \clock_counter[0]_net_1 ), .Y(N_144));
    CLKINT output_signal_RNI2QGD (.A(output_signal_0), .Y(
        output_signal_c));
    OR3A \clock_counter_RNI3U8B[5]  (.A(\clock_counter[5]_net_1 ), .B(
        N_42), .C(N_45), .Y(N_46));
    XAI1 \counter_RNO_0[1]  (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(trigger_signal_c), .Y(counter_n1_i_0));
    AOI1 \counter_RNO[1]  (.A(N_123_1), .B(N_151), .C(counter_n1_i_0), 
        .Y(N_5));
    DFN1E1C0 \clock_counter[9]  (.D(clock_counter_n9), .CLK(
        ref_signal_c), .CLR(reset_c), .E(clock_countere), .Q(
        \clock_counter[9]_net_1 ));
    DFN1E1C0 \clock_counter[15]  (.D(clock_counter_n15), .CLK(
        ref_signal_c), .CLR(reset_c), .E(clock_countere), .Q(
        \clock_counter[15]_net_1 ));
    XA1A \clock_counter_RNO[12]  (.A(un6lto12), .B(N_49), .C(
        trigger_signal_c), .Y(clock_counter_n12));
    XA1A \clock_counter_RNO[13]  (.A(\clock_counter[13]_net_1 ), .B(
        N_50), .C(trigger_signal_c), .Y(clock_counter_n13));
    AO1B \counter_RNISQHA3[0]  (.A(counter_0_sqmuxa_i_a2_0), .B(N_151), 
        .C(trigger_signal_c), .Y(N_8));
    OA1 output_signal_RNO_2 (.A(N_45), .B(N_150), .C(
        output_signal_1_sqmuxa_i_a2_2), .Y(N_145));
    XA1A \clock_counter_RNO[14]  (.A(\clock_counter[14]_net_1 ), .B(
        N_52), .C(trigger_signal_c), .Y(clock_counter_n14));
    DFN1E1C0 \clock_counter[5]  (.D(N_23), .CLK(ref_signal_c), .CLR(
        reset_c), .E(clock_countere), .Q(\clock_counter[5]_net_1 ));
    OR2A output_signal_RNO_10 (.A(trigger_signal_c), .B(
        \clock_counter[13]_net_1 ), .Y(N_36_3));
    OR3 output_signal_RNO_4 (.A(\clock_counter[14]_net_1 ), .B(
        \clock_counter[15]_net_1 ), .C(N_36_3), .Y(
        output_signal_1_sqmuxa_i_1));
    XA1A \clock_counter_RNO[5]  (.A(\clock_counter[5]_net_1 ), .B(N_42)
        , .C(counter_n0), .Y(N_23));
    OR2 \clock_counter_RNIFVF2_0[1]  (.A(\clock_counter[1]_net_1 ), .B(
        \clock_counter[0]_net_1 ), .Y(N_51));
    NOR2B \counter_RNI1ROV[5]  (.A(\counter[5]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(N_123_1));
    OR2A \clock_counter_RNO_0[15]  (.A(\clock_counter[14]_net_1 ), .B(
        N_52), .Y(N_91));
    NOR2 output_signal_RNO_12 (.A(\clock_counter[4]_net_1 ), .B(
        \clock_counter[5]_net_1 ), .Y(output_signal_1_sqmuxa_i_a2_3_0));
    DFN1C0 \counter[4]  (.D(counter_n4), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[4]_net_1 ));
    DFN1C0 \counter[5]  (.D(counter_n5), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[5]_net_1 ));
    XA1A \clock_counter_RNO[10]  (.A(\clock_counter[10]_net_1 ), .B(
        N_61), .C(trigger_signal_c), .Y(clock_counter_n10));
    XA1B \counter_RNO[2]  (.A(counter_c1), .B(\counter[2]_net_1 ), .C(
        N_8), .Y(counter_n2));
    OR2 \clock_counter_RNIB3OL[10]  (.A(N_47), .B(N_46), .Y(N_48));
    NOR2B output_signal_RNO_5 (.A(un6lto11), .B(un6lto12), .Y(N_147));
    NOR3 output_signal_RNO (.A(N_146), .B(output_signal_1_sqmuxa_i_3), 
        .C(N_145), .Y(N_36));
    GND GND_i (.Y(GND));
    XA1B \counter_RNO[5]  (.A(counter_44_0), .B(\counter[5]_net_1 ), 
        .C(N_8), .Y(counter_n5));
    XA1B \counter_RNO[3]  (.A(counter_c2), .B(\counter[3]_net_1 ), .C(
        N_8), .Y(counter_n3));
    NOR2B \counter_RNIPIOV[1]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(counter_c1));
    OR2A \clock_counter_RNO_0[10]  (.A(\clock_counter[9]_net_1 ), .B(
        N_46), .Y(N_61));
    OR2B \clock_counter_RNIFVF2[1]  (.A(\clock_counter[1]_net_1 ), .B(
        \clock_counter[0]_net_1 ), .Y(N_39));
    NOR2B output_signal_RNO_11 (.A(\clock_counter[8]_net_1 ), .B(
        un6lto7), .Y(output_signal_1_sqmuxa_i_a2_2_0));
    DFN1C0 \counter[1]  (.D(N_5), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[1]_net_1 ));
    XA1A \clock_counter_RNO[3]  (.A(\clock_counter[3]_net_1 ), .B(N_40)
        , .C(counter_n0), .Y(N_27));
    DFN1E1C0 \clock_counter[2]  (.D(N_29), .CLK(ref_signal_c), .CLR(
        reset_c), .E(clock_countere), .Q(\clock_counter[2]_net_1 ));
    OR3 output_signal_RNO_1 (.A(output_signal_1_sqmuxa_i_1), .B(N_147), 
        .C(N_148), .Y(output_signal_1_sqmuxa_i_3));
    NOR2B \counter_RNO_0[5]  (.A(\counter[4]_net_1 ), .B(counter_c3), 
        .Y(counter_44_0));
    DFN1C0 \counter[3]  (.D(counter_n3), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[3]_net_1 ));
    AO1B \counter_RNISQHA3[5]  (.A(clock_counterlde_0_a2_1), .B(N_151), 
        .C(trigger_signal_c), .Y(clock_countere));
    NOR3 \counter_RNIQ0LF1[1]  (.A(\counter[2]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[1]_net_1 ), .Y(N_151));
    DFN1E1C0 \clock_counter[7]  (.D(N_19), .CLK(ref_signal_c), .CLR(
        reset_c), .E(clock_countere), .Q(un6lto7));
    DFN1E1C0 \clock_counter[14]  (.D(clock_counter_n14), .CLK(
        ref_signal_c), .CLR(reset_c), .E(clock_countere), .Q(
        \clock_counter[14]_net_1 ));
    XA1A \clock_counter_RNO[7]  (.A(un6lto7), .B(N_53), .C(counter_n0), 
        .Y(N_19));
    OR2 \clock_counter_RNI2305[1]  (.A(output_signal_1_sqmuxa_i_o2_0), 
        .B(N_51), .Y(N_55));
    NOR3A output_signal_RNO_8 (.A(output_signal_1_sqmuxa_i_a2_1), .B(
        \clock_counter[9]_net_1 ), .C(\clock_counter[10]_net_1 ), .Y(
        output_signal_1_sqmuxa_i_a2_2));
    NOR2B \counter_RNIT3LF1[0]  (.A(\counter[0]_net_1 ), .B(N_123_1), 
        .Y(counter_0_sqmuxa_i_a2_0));
    OA1C \clock_counter_RNO_0[8]  (.A(un6lto7), .B(N_53), .C(
        \clock_counter[8]_net_1 ), .Y(N_137));
    OR2A \clock_counter_RNIO0O3[2]  (.A(\clock_counter[2]_net_1 ), .B(
        N_39), .Y(N_40));
    OR3C \clock_counter_RNIAJO3[6]  (.A(\clock_counter[8]_net_1 ), .B(
        \clock_counter[6]_net_1 ), .C(un6lto7), .Y(N_45));
    DFN1E1C0 \clock_counter[12]  (.D(clock_counter_n12), .CLK(
        ref_signal_c), .CLR(reset_c), .E(clock_countere), .Q(un6lto12));
    NOR3B output_signal_RNO_0 (.A(N_55), .B(
        output_signal_1_sqmuxa_i_a2_0_2), .C(N_47), .Y(N_146));
    NOR3B \clock_counter_RNO[8]  (.A(N_46), .B(counter_n0), .C(N_137), 
        .Y(N_17));
    NOR3C output_signal_RNO_9 (.A(\clock_counter[5]_net_1 ), .B(
        \clock_counter[4]_net_1 ), .C(un6lto12), .Y(
        output_signal_1_sqmuxa_i_a2_0_1));
    DFN1E1C0 output_signal (.D(N_36), .CLK(ref_signal_c), .CLR(reset_c)
        , .E(clock_countere), .Q(output_signal_0));
    OR2A \clock_counter_RNIUV581[12]  (.A(un6lto12), .B(N_49), .Y(N_50)
        );
    DFN1E1C0 \clock_counter[13]  (.D(clock_counter_n13), .CLK(
        ref_signal_c), .CLR(reset_c), .E(clock_countere), .Q(
        \clock_counter[13]_net_1 ));
    XA1A \clock_counter_RNO[9]  (.A(\clock_counter[9]_net_1 ), .B(N_46)
        , .C(trigger_signal_c), .Y(clock_counter_n9));
    XA1A \clock_counter_RNO[11]  (.A(un6lto11), .B(N_48), .C(
        trigger_signal_c), .Y(clock_counter_n11));
    DFN1E1C0 \clock_counter[11]  (.D(clock_counter_n11), .CLK(
        ref_signal_c), .CLR(reset_c), .E(clock_countere), .Q(un6lto11));
    NOR3C output_signal_RNO_3 (.A(\clock_counter[8]_net_1 ), .B(
        \clock_counter[6]_net_1 ), .C(output_signal_1_sqmuxa_i_a2_0_1), 
        .Y(output_signal_1_sqmuxa_i_a2_0_2));
    OA1C \clock_counter_RNO_0[6]  (.A(\clock_counter[5]_net_1 ), .B(
        N_42), .C(\clock_counter[6]_net_1 ), .Y(N_139));
    XA1 \clock_counter_RNO[1]  (.A(\clock_counter[0]_net_1 ), .B(
        \clock_counter[1]_net_1 ), .C(counter_n0), .Y(N_31));
    OR2A \clock_counter_RNIPVCH1[13]  (.A(\clock_counter[13]_net_1 ), 
        .B(N_50), .Y(N_52));
    NOR2A \counter_RNI1V3R[0]  (.A(trigger_signal_c), .B(
        \counter[0]_net_1 ), .Y(counter_n0));
    NOR3B output_signal_RNO_6 (.A(output_signal_1_sqmuxa_i_a2_2_0), .B(
        un6lto12), .C(N_47), .Y(N_148));
    XA1A \clock_counter_RNO[15]  (.A(\clock_counter[15]_net_1 ), .B(
        N_91), .C(trigger_signal_c), .Y(clock_counter_n15));
    DFN1E1C0 \clock_counter[10]  (.D(clock_counter_n10), .CLK(
        ref_signal_c), .CLR(reset_c), .E(clock_countere), .Q(
        \clock_counter[10]_net_1 ));
    XA1A \clock_counter_RNO[2]  (.A(\clock_counter[2]_net_1 ), .B(N_39)
        , .C(counter_n0), .Y(N_29));
    NOR2B \counter_RNIM9HV1[3]  (.A(counter_c2), .B(\counter[3]_net_1 )
        , .Y(counter_c3));
    DFN1C0 \counter[0]  (.D(counter_n0), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[0]_net_1 ));
    NOR3B \clock_counter_RNO[6]  (.A(counter_n0), .B(N_53), .C(N_139), 
        .Y(N_21));
    NOR2 output_signal_RNO_13 (.A(un6lto11), .B(un6lto12), .Y(
        output_signal_1_sqmuxa_i_a2_1));
    OR2B \clock_counter_RNI85FA[10]  (.A(\clock_counter[10]_net_1 ), 
        .B(\clock_counter[9]_net_1 ), .Y(N_47));
    
endmodule


module demodulator(
       demodulator_0_ord,
       demodulator_0_ctg,
       demodulator_0_cur_flag,
       demodulator_0_cur_scheme,
       reset_c,
       ref_signal_c,
       insig_c,
       mac_0_working
    );
output [1:0] demodulator_0_ord;
output [1:0] demodulator_0_ctg;
output [7:0] demodulator_0_cur_flag;
output [47:0] demodulator_0_cur_scheme;
input  reset_c;
input  ref_signal_c;
input  insig_c;
input  mac_0_working;

    wire un1_working_2_1, un1_buffer22, un1_working_2_0, 
        un1_counter11_1_0, buffer_3_sqmuxa_2, len_3_sqmuxa_1_0, 
        un1_counter11_0, un1_counter11_0_0, cur_scheme_1_sqmuxa_0, 
        cur_scheme_0_sqmuxa, counter10, \DWACT_ADD_CI_0_g_array_2[0] , 
        \DWACT_ADD_CI_0_g_array_1[0] , \DWACT_ADD_CI_0_pog_array_1[0] , 
        \DWACT_ADD_CI_0_TMP[0] , \len[1]_net_1 , 
        \DWACT_ADD_CI_0_g_array_12[0] , \len[2]_net_1 , 
        \DWACT_ADD_CI_0_g_array_12_1[0] , \len[4]_net_1 , N_5, 
        \counter[1]_net_1 , \counter[0]_net_1 , N_3, 
        \counter[3]_net_1 , \DWACT_FINC_E[0] , cur_flag_1_sqmuxa_i, 
        cur_flag_1_sqmuxa, ord_1_sqmuxa_0, un1_insig_i_0, 
        waittimelde_i_o2_1, ord36, ord35, ord34, checksum_4_iv_0_0, 
        checksum_4_iv_0_a4_1_0, buffer22, N_76, latency_n5_i_0, 
        \latency[5]_net_1 , N_42, latency_n1_i_0, \latency[0]_net_1 , 
        \latency[1]_net_1 , latency_n4_i_0, N_40, \latency[3]_net_1 , 
        \latency[4]_net_1 , latency_n3_i_0, latency_n2_i_0, 
        \latency[2]_net_1 , N_56, checksum_net_1, 
        cur_scheme_0_sqmuxa_1, \buffer[49]_net_1 , \buffer[50]_net_1 , 
        un1_LOWERBOUND_0_1_3, un1_LOWERBOUND_0_1_2, N_48, 
        un1_LOWERBOUND_0lto9_2, un1_LOWERBOUND_0lto9_5, 
        un1_LOWERBOUND_0lto9_4, counter10_2, counter10_1, 
        \counter[2]_net_1 , counter10_0, \counter[5]_net_1 , 
        \counter[4]_net_1 , cur_flag_0_sqmuxa_1, \buffer[10]_net_1 , 
        \buffer[9]_net_1 , un1_buffer21_3_i_i_o2_5, 
        un1_buffer21_3_i_i_o2_1, un1_buffer21_3_i_i_o2_0, 
        un1_buffer21_3_i_i_o2_4, \latency[9]_net_1 , 
        \latency[6]_net_1 , N_39, \latency[8]_net_1 , 
        \latency[7]_net_1 , buffer21_8, buffer21_2, buffer21_1, 
        buffer21_5, buffer21_7, \waittime[4]_net_1 , buffer21_4, 
        \waittime[9]_net_1 , \waittime[7]_net_1 , \waittime[6]_net_1 , 
        \waittime[10]_net_1 , \waittime[5]_net_1 , \waittime[2]_net_1 , 
        \waittime[1]_net_1 , \waittime[3]_net_1 , \waittime[8]_net_1 , 
        \waittime[0]_net_1 , ord36_0_a2_0, \len[5]_net_1 , 
        un1_LOWERBOUND_0lt9_1, un1_LOWERBOUND_0lt9_0, ord35_0_a2_0, 
        \len[3]_net_1 , N_18, ord10, \buffer[1]_net_1 , 
        \buffer[2]_net_1 , N_61, N_79, buffer21, N_16, 
        cur_flag_0_sqmuxa, \len[0]_net_1 , ord_1_sqmuxa, 
        un1_cur_scheme_0_sqmuxa, N_13, len_3_sqmuxa, len_3_sqmuxa_1, 
        N_75_1, cur_scheme_1_sqmuxa, ctg_0_sqmuxa, 
        \len_RNI2H48I[3]_net_1 , un1_counter11, checksum_4, N_58_i, 
        un1_LOWERBOUND_0lto9, N_19, N_54, N_278, N_21, N_44, N_23, 
        N_43, N_25, N_27, N_29, N_31, N_33, waittime_n2, waittime_c1, 
        latency_1_sqmuxa_1, waittime_n3, waittime_c2, waittime_n4, 
        waittime_c3, waittime_n5, waittime_c4, waittime_n6, 
        waittime_c5, waittime_n7, waittime_c6, waittime_n8, 
        waittime_c7, waittime_n9, waittime_c8, waittime_n10, 
        waittime_22_0, \buffer_9[4] , \buffer[3]_net_1 , \buffer_9[8] , 
        \buffer[7]_net_1 , \buffer_9[12] , \buffer[11]_net_1 , 
        \buffer_9[13] , \buffer[12]_net_1 , \buffer_9[14] , 
        \buffer[13]_net_1 , \buffer_9[15] , \buffer[14]_net_1 , 
        \buffer_9[16] , \buffer[15]_net_1 , \buffer_9[17] , 
        \buffer[16]_net_1 , \buffer_9[18] , \buffer[17]_net_1 , 
        \buffer_9[19] , \buffer[18]_net_1 , \buffer_9[20] , 
        \buffer[19]_net_1 , \buffer_9[21] , \buffer[20]_net_1 , 
        \buffer_9[22] , \buffer[21]_net_1 , \buffer_9[23] , 
        \buffer[22]_net_1 , \buffer_9[24] , \buffer[23]_net_1 , 
        \buffer_9[25] , \buffer[24]_net_1 , \buffer_9[26] , 
        \buffer[25]_net_1 , \buffer_9[27] , \buffer[26]_net_1 , 
        \buffer_9[28] , \buffer[27]_net_1 , \buffer_9[29] , 
        \buffer[28]_net_1 , \buffer_9[30] , \buffer[29]_net_1 , 
        \buffer_9[31] , \buffer[30]_net_1 , \buffer_9[32] , 
        \buffer[31]_net_1 , \buffer_9[33] , \buffer[32]_net_1 , 
        \buffer_9[34] , \buffer[33]_net_1 , \buffer_9[35] , 
        \buffer[34]_net_1 , un1_working_2, \buffer_9[36] , 
        \buffer[35]_net_1 , \buffer_9[37] , \buffer[36]_net_1 , 
        \buffer_9[38] , \buffer[37]_net_1 , \buffer_9[39] , 
        \buffer[38]_net_1 , \buffer_9[40] , \buffer[39]_net_1 , 
        \buffer_9[41] , \buffer[40]_net_1 , \buffer_9[42] , 
        \buffer[41]_net_1 , \buffer_9[43] , \buffer[42]_net_1 , 
        \buffer_9[44] , \buffer[43]_net_1 , \buffer_9[45] , 
        \buffer[44]_net_1 , \buffer_9[46] , \buffer[45]_net_1 , 
        \buffer_9[47] , \buffer[46]_net_1 , \buffer_9[48] , 
        \buffer[47]_net_1 , \buffer_9[49] , \buffer[48]_net_1 , 
        \buffer_9[3] , \buffer_9[10] , \buffer_9[11] , \buffer_9[50] , 
        \buffer_9[1] , \buffer[0]_net_1 , \buffer_9[7] , 
        \buffer[6]_net_1 , \buffer_9[6] , \buffer[5]_net_1 , N_577, 
        waittime_n1, \buffer_9[9] , \buffer[8]_net_1 , N_37, N_8, 
        checksum_2_sqmuxa, latency_n9, N_55, \len_10[2] , I_23, 
        un1_len_1_sqmuxa, \len_10[3] , I_22, \len_10[4] , I_21, 
        \len_10[5] , I_26, \counter_3[1] , I_5, \counter_3[4] , I_12, 
        \counter_3[5] , I_14, \len_10[0] , 
        \DWACT_ADD_CI_0_partial_sum[0] , \len_10[1] , I_24, 
        un1_buffer21_1, checksum_0_sqmuxa, \buffer_9[2] , N_73, 
        \buffer_9[5] , \buffer[4]_net_1 , I_4, I_7, I_9, 
        \DWACT_ADD_CI_0_partial_sum_0[0] , \ord_11[1] , 
        \DWACT_ADD_CI_0_TMP_0[0] , N_2, N_4, GND, VCC;
    
    NOR2A \buffer_RNO[49]  (.A(\buffer[48]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[49] ));
    DFN1E0C0 \latency[7]  (.D(N_21), .CLK(ref_signal_c), .CLR(reset_c), 
        .E(N_8), .Q(\latency[7]_net_1 ));
    NOR2A \buffer_RNO[3]  (.A(\buffer[2]_net_1 ), .B(un1_working_2_0), 
        .Y(\buffer_9[3] ));
    NOR3C \waittime_RNI9V1F1[1]  (.A(buffer21_2), .B(buffer21_1), .C(
        buffer21_5), .Y(buffer21_8));
    DFN1E0C0 \buffer[24]  (.D(\buffer_9[24] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[24]_net_1 ));
    NOR2A \buffer_RNO[17]  (.A(\buffer[16]_net_1 ), .B(un1_working_2_0)
        , .Y(\buffer_9[17] ));
    OR2A \latency_RNICS5DM[9]  (.A(un1_buffer22), .B(mac_0_working), 
        .Y(un1_working_2));
    DFN1E1C0 checksum (.D(checksum_4), .CLK(ref_signal_c), .CLR(
        reset_c), .E(counter10), .Q(checksum_net_1));
    XA1 \waittime_RNO[5]  (.A(waittime_c4), .B(\waittime[5]_net_1 ), 
        .C(latency_1_sqmuxa_1), .Y(waittime_n5));
    DFN1E0C0 \buffer[3]  (.D(\buffer_9[3] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(un1_counter11_0_0), .Q(\buffer[3]_net_1 ));
    AND2 ord_11_I_1 (.A(demodulator_0_ord[0]), .B(ord_1_sqmuxa), .Y(
        \DWACT_ADD_CI_0_TMP_0[0] ));
    NOR2A \buffer_RNO[9]  (.A(\buffer[8]_net_1 ), .B(un1_working_2_0), 
        .Y(\buffer_9[9] ));
    DFN1C0 \len[4]  (.D(\len_10[4] ), .CLK(ref_signal_c), .CLR(reset_c)
        , .Q(\len[4]_net_1 ));
    OR2A \latency_RNICS5DM_0[9]  (.A(un1_buffer22), .B(mac_0_working), 
        .Y(un1_working_2_1));
    NOR2A \buffer_RNO[35]  (.A(\buffer[34]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[35] ));
    DFN1E0C0 \buffer[41]  (.D(\buffer_9[41] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[41]_net_1 ));
    DFN1E0C0 \latency[8]  (.D(N_19), .CLK(ref_signal_c), .CLR(reset_c), 
        .E(N_8), .Q(\latency[8]_net_1 ));
    DFN1E1C0 \cur_scheme[43]  (.D(\buffer[44]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[43]));
    NOR2A \buffer_RNO[25]  (.A(\buffer[24]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[25] ));
    DFN1E1C0 \cur_scheme[41]  (.D(\buffer[42]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[41]));
    DFN1E0C0 \buffer[10]  (.D(\buffer_9[10] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_0_0), .Q(\buffer[10]_net_1 ));
    DFN1E0C0 \latency[3]  (.D(N_29), .CLK(ref_signal_c), .CLR(reset_c), 
        .E(N_8), .Q(\latency[3]_net_1 ));
    DFN1E0C0 \buffer[9]  (.D(\buffer_9[9] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(un1_counter11_0_0), .Q(\buffer[9]_net_1 ));
    NOR2A \buffer_RNO[47]  (.A(\buffer[46]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[47] ));
    DFN1E0C0 \buffer[43]  (.D(\buffer_9[43] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[43]_net_1 ));
    NOR3B \len_RNIFUSA[0]  (.A(\len[1]_net_1 ), .B(\len[0]_net_1 ), .C(
        \len[2]_net_1 ), .Y(N_16));
    DFN1E0C0 \buffer[31]  (.D(\buffer_9[31] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[31]_net_1 ));
    INV un3_counter_I_4 (.A(\counter[0]_net_1 ), .Y(I_4));
    DFN1E1C0 \cur_scheme[7]  (.D(\buffer[8]_net_1 ), .CLK(ref_signal_c)
        , .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[7]));
    DFN1E1C0 \cur_scheme[46]  (.D(\buffer[47]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[46]));
    NOR2B \buffer_RNIFLVF1[9]  (.A(cur_flag_0_sqmuxa_1), .B(ord35), .Y(
        cur_flag_0_sqmuxa));
    AND3 un3_counter_I_10 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(
        \DWACT_FINC_E[0] ));
    DFN1E1C0 \cur_scheme[6]  (.D(\buffer[7]_net_1 ), .CLK(ref_signal_c)
        , .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[6]));
    DFN1E0C0 \buffer[33]  (.D(\buffer_9[33] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[33]_net_1 ));
    DFN1E1C0 \cur_scheme[4]  (.D(\buffer[5]_net_1 ), .CLK(ref_signal_c)
        , .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[4]));
    NOR2 \buffer_RNIME533[9]  (.A(cur_scheme_0_sqmuxa), .B(
        cur_flag_0_sqmuxa), .Y(buffer_3_sqmuxa_2));
    DFN1E0C0 \buffer[45]  (.D(\buffer_9[45] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[45]_net_1 ));
    NOR2B \len_RNIHR87[5]  (.A(\len[5]_net_1 ), .B(\len[4]_net_1 ), .Y(
        ord36_0_a2_0));
    XA1 \waittime_RNO[9]  (.A(waittime_c8), .B(\waittime[9]_net_1 ), 
        .C(latency_1_sqmuxa_1), .Y(waittime_n9));
    NOR2A \waittime_RNIU8NJ2[4]  (.A(un1_insig_i_0), .B(buffer21), .Y(
        latency_1_sqmuxa_1));
    DFN1E1C0 \cur_scheme[25]  (.D(\buffer[26]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[25]));
    DFN1E0C0 \buffer[35]  (.D(\buffer_9[35] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[35]_net_1 ));
    XOR2 un1_len_1_I_23 (.A(\len[2]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_1[0] ), .Y(I_23));
    AND3 un3_counter_I_13 (.A(\DWACT_FINC_E[0] ), .B(
        \counter[3]_net_1 ), .C(\counter[4]_net_1 ), .Y(N_2));
    NOR2A \buffer_RNO[50]  (.A(\buffer[49]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[50] ));
    NOR2A \counter_RNIBJ18[1]  (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .Y(counter10_2));
    DFN1E0C0 \buffer[16]  (.D(\buffer_9[16] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_0_0), .Q(\buffer[16]_net_1 ));
    DFN1E1C0 \cur_scheme[8]  (.D(\buffer[9]_net_1 ), .CLK(ref_signal_c)
        , .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[8]));
    DFN1C0 \counter[3]  (.D(I_9), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[3]_net_1 ));
    DFN1C0 \counter[2]  (.D(I_7), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[2]_net_1 ));
    AO1D \latency_RNIUD5OC_0[9]  (.A(un1_buffer21_3_i_i_o2_5), .B(
        un1_buffer21_3_i_i_o2_4), .C(un1_buffer21_1), .Y(N_13));
    NOR3B \len_RNI76QL[3]  (.A(N_16), .B(N_18), .C(\len[3]_net_1 ), .Y(
        ord34));
    NOR3C \buffer_RNINDNFF[9]  (.A(cur_flag_0_sqmuxa), .B(counter10), 
        .C(len_3_sqmuxa_1_0), .Y(cur_flag_1_sqmuxa));
    NOR2B \len_RNO[3]  (.A(I_22), .B(un1_len_1_sqmuxa), .Y(\len_10[3] )
        );
    NOR2A \buffer_RNO[34]  (.A(\buffer[33]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[34] ));
    DFN1E0C0 \buffer[18]  (.D(\buffer_9[18] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[18]_net_1 ));
    DFN1E1C0 \cur_scheme[19]  (.D(\buffer[20]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[19]));
    NOR2B un1_len_1_I_29 (.A(\DWACT_ADD_CI_0_g_array_2[0] ), .B(
        \len[4]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12_1[0] ));
    NOR2A \buffer_RNO[24]  (.A(\buffer[23]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[24] ));
    NOR2A \buffer_RNO[4]  (.A(\buffer[3]_net_1 ), .B(un1_working_2_0), 
        .Y(\buffer_9[4] ));
    DFN1E0C0 \buffer[27]  (.D(\buffer_9[27] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[27]_net_1 ));
    DFN1E0C0 \waittime[5]  (.D(waittime_n5), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_37), .Q(\waittime[5]_net_1 ));
    DFN1E1C0 \cur_scheme[20]  (.D(\buffer[21]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[20]));
    AO1C \counter_RNIAAI71[1]  (.A(mac_0_working), .B(insig_c), .C(
        counter10), .Y(un1_counter11_0));
    AO1 \counter_RNIRAAIH_0[1]  (.A(buffer_3_sqmuxa_2), .B(
        len_3_sqmuxa_1_0), .C(un1_counter11_0), .Y(un1_counter11_1_0));
    NOR2A \waittime_RNIF5J52[4]  (.A(buffer21), .B(insig_c), .Y(
        checksum_0_sqmuxa));
    NOR2A \buffer_RNO[8]  (.A(\buffer[7]_net_1 ), .B(un1_working_2_0), 
        .Y(\buffer_9[8] ));
    XA1 \waittime_RNO[4]  (.A(waittime_c3), .B(\waittime[4]_net_1 ), 
        .C(latency_1_sqmuxa_1), .Y(waittime_n4));
    XA1 \waittime_RNO[10]  (.A(waittime_22_0), .B(\waittime[10]_net_1 )
        , .C(latency_1_sqmuxa_1), .Y(waittime_n10));
    XOR2 un3_counter_I_14 (.A(N_2), .B(\counter[5]_net_1 ), .Y(I_14));
    NOR2A \buffer_RNO[30]  (.A(\buffer[29]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[30] ));
    NOR2A \counter_RNO[1]  (.A(I_5), .B(counter10), .Y(\counter_3[1] ));
    NOR2A \buffer_RNO[20]  (.A(\buffer[19]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[20] ));
    DFN1C0 \counter[4]  (.D(\counter_3[4] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[4]_net_1 ));
    XOR2 un3_counter_I_5 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .Y(I_5));
    DFN1E1C0 \cur_scheme[27]  (.D(\buffer[28]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[27]));
    OR2A \counter_RNIBFSB3[1]  (.A(counter10), .B(latency_1_sqmuxa_1), 
        .Y(N_8));
    NOR2B \waittime_RNI4VFA1[7]  (.A(waittime_c6), .B(
        \waittime[7]_net_1 ), .Y(waittime_c7));
    DFN1E1C0 \cur_scheme[35]  (.D(\buffer[36]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[35]));
    DFN1E0C0 \buffer[40]  (.D(\buffer_9[40] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[40]_net_1 ));
    DFN1E0C0 \buffer[14]  (.D(\buffer_9[14] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_0_0), .Q(\buffer[14]_net_1 ));
    NOR2A \buffer_RNO[5]  (.A(\buffer[4]_net_1 ), .B(un1_working_2_0), 
        .Y(\buffer_9[5] ));
    NOR2 \latency_RNO[4]  (.A(latency_n4_i_0), .B(N_278), .Y(N_27));
    GND GND_i (.Y(GND));
    DFN1E1C0 \cur_scheme[12]  (.D(\buffer[13]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[12]));
    XA1 \waittime_RNO[8]  (.A(waittime_c7), .B(\waittime[8]_net_1 ), 
        .C(latency_1_sqmuxa_1), .Y(waittime_n8));
    AND2 un1_len_1_I_1 (.A(\len[0]_net_1 ), .B(\len_RNI2H48I[3]_net_1 )
        , .Y(\DWACT_ADD_CI_0_TMP[0] ));
    DFN1E0C0 \buffer[30]  (.D(\buffer_9[30] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[30]_net_1 ));
    DFN1E1C0 \cur_scheme[5]  (.D(\buffer[6]_net_1 ), .CLK(ref_signal_c)
        , .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[5]));
    DFN1E1C0 \cur_scheme[14]  (.D(\buffer[15]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[14]));
    NOR2B \waittime_RNIJPJA[1]  (.A(\waittime[0]_net_1 ), .B(
        \waittime[1]_net_1 ), .Y(waittime_c1));
    NOR2B checksum_RNO_2 (.A(checksum_net_1), .B(un1_insig_i_0), .Y(
        checksum_4_iv_0_a4_1_0));
    DFN1E1C0 \cur_flag[7]  (.D(\buffer[8]_net_1 ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(cur_flag_1_sqmuxa), .Q(
        demodulator_0_cur_flag[7]));
    OR2B \latency_RNIBOKM[0]  (.A(\latency[1]_net_1 ), .B(
        \latency[0]_net_1 ), .Y(N_56));
    XOR2 ord_11_I_10 (.A(demodulator_0_ord[1]), .B(
        \DWACT_ADD_CI_0_TMP_0[0] ), .Y(\ord_11[1] ));
    DFN1E1C0 \cur_scheme[30]  (.D(\buffer[31]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[30]));
    NOR2B \counter_RNIAAI71_0[1]  (.A(un1_insig_i_0), .B(counter10), 
        .Y(ord_1_sqmuxa_0));
    NOR2A \buffer_RNO[0]  (.A(N_79), .B(mac_0_working), .Y(
        checksum_2_sqmuxa));
    DFN1C0 \len[0]  (.D(\len_10[0] ), .CLK(ref_signal_c), .CLR(reset_c)
        , .Q(\len[0]_net_1 ));
    DFN1E0C0 \latency[9]  (.D(latency_n9), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_8), .Q(\latency[9]_net_1 ));
    NOR2B un3_counter_I_6 (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(N_5));
    DFN1E1C0 \cur_scheme[18]  (.D(\buffer[19]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[18]));
    NOR3 \latency_RNIUD5OC[9]  (.A(un1_buffer21_3_i_i_o2_4), .B(
        un1_buffer21_3_i_i_o2_5), .C(un1_buffer21_1), .Y(N_79));
    NOR2A \buffer_RNO[18]  (.A(\buffer[17]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[18] ));
    DFN1E1C0 \cur_scheme[23]  (.D(\buffer[24]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[23]));
    DFN1E0C0 \latency[6]  (.D(N_23), .CLK(ref_signal_c), .CLR(reset_c), 
        .E(N_8), .Q(\latency[6]_net_1 ));
    DFN1E1C0 \cur_scheme[21]  (.D(\buffer[22]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[21]));
    AX1D checksum_RNO_0 (.A(un1_buffer21_3_i_i_o2_4), .B(
        un1_buffer21_3_i_i_o2_5), .C(checksum_net_1), .Y(N_58_i));
    DFN1E0C0 \buffer[29]  (.D(\buffer_9[29] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[29]_net_1 ));
    DFN1E1C0 \cur_scheme[37]  (.D(\buffer[38]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[37]));
    AND3 un3_counter_I_8 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(N_4));
    DFN1E0C0 \buffer[46]  (.D(\buffer_9[46] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[46]_net_1 ));
    DFN1E0C0 \waittime[1]  (.D(waittime_n1), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_37), .Q(\waittime[1]_net_1 ));
    NOR2A \buffer_RNO[48]  (.A(\buffer[47]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[48] ));
    NOR2A \buffer_RNO[2]  (.A(\buffer[1]_net_1 ), .B(un1_working_2_0), 
        .Y(\buffer_9[2] ));
    OR2 \latency_RNIR8LM[9]  (.A(\latency[8]_net_1 ), .B(
        \latency[9]_net_1 ), .Y(un1_LOWERBOUND_0lto9_5));
    DFN1E0C0 \waittime[2]  (.D(waittime_n2), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_37), .Q(\waittime[2]_net_1 ));
    NOR3B \len_RNI76QL_0[3]  (.A(N_16), .B(ord36_0_a2_0), .C(
        \len[3]_net_1 ), .Y(ord36));
    DFN1E0C0 \waittime[7]  (.D(waittime_n7), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_37), .Q(\waittime[7]_net_1 ));
    NOR2A \buffer_RNO[11]  (.A(\buffer[10]_net_1 ), .B(un1_working_2_0)
        , .Y(\buffer_9[11] ));
    DFN1E0C0 \buffer[5]  (.D(\buffer_9[5] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(un1_counter11_0_0), .Q(\buffer[5]_net_1 ));
    DFN1E1C0 \cur_scheme[26]  (.D(\buffer[27]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[26]));
    NOR2A \buffer_RNO[39]  (.A(\buffer[38]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[39] ));
    NOR2A \buffer_RNO[1]  (.A(\buffer[0]_net_1 ), .B(un1_working_2_0), 
        .Y(\buffer_9[1] ));
    DFN1E0C0 \buffer[50]  (.D(\buffer_9[50] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[50]_net_1 ));
    NOR2A \buffer_RNO[29]  (.A(\buffer[28]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[29] ));
    DFN1E0C0 \buffer[48]  (.D(\buffer_9[48] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[48]_net_1 ));
    OR2A \latency_RNO_0[9]  (.A(\latency[8]_net_1 ), .B(N_54), .Y(N_55)
        );
    NOR3B \latency_RNIVAS69[0]  (.A(un1_LOWERBOUND_0lto9), .B(
        un1_LOWERBOUND_0_1_3), .C(buffer21), .Y(buffer22));
    VCC VCC_i (.Y(VCC));
    DFN1E0C0 \buffer[36]  (.D(\buffer_9[36] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[36]_net_1 ));
    NOR2B \waittime_RNIL3QF1[8]  (.A(waittime_c7), .B(
        \waittime[8]_net_1 ), .Y(waittime_c8));
    OR2A \latency_RNI4QJQ2[7]  (.A(\latency[7]_net_1 ), .B(N_44), .Y(
        N_54));
    DFN1C0 \counter[1]  (.D(\counter_3[1] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[1]_net_1 ));
    NOR2 \waittime_RNIMSJA[1]  (.A(\waittime[1]_net_1 ), .B(
        \waittime[3]_net_1 ), .Y(buffer21_2));
    OR2 \latency_RNITO1VL[9]  (.A(buffer22), .B(N_79), .Y(un1_buffer22)
        );
    NOR3A \latency_RNIV29H3[2]  (.A(un1_LOWERBOUND_0_1_2), .B(N_48), 
        .C(un1_LOWERBOUND_0lto9_2), .Y(un1_LOWERBOUND_0_1_3));
    DFN1E1C0 \cur_scheme[3]  (.D(\buffer[4]_net_1 ), .CLK(ref_signal_c)
        , .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[3]));
    NOR2A \counter_RNO[5]  (.A(I_14), .B(counter10), .Y(\counter_3[5] )
        );
    NOR2A \buffer_RNO[41]  (.A(\buffer[40]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[41] ));
    OR2A \latency_RNI26V11[1]  (.A(\latency[1]_net_1 ), .B(N_39), .Y(
        N_40));
    DFN1E0C0 \buffer[38]  (.D(\buffer_9[38] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[38]_net_1 ));
    NOR2B un1_len_1_I_27 (.A(\DWACT_ADD_CI_0_TMP[0] ), .B(
        \len[1]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_1[0] ));
    NOR3B \waittime_RNIP1QP[10]  (.A(\waittime[7]_net_1 ), .B(
        \waittime[6]_net_1 ), .C(\waittime[10]_net_1 ), .Y(buffer21_5));
    DFN1E0C0 \buffer[17]  (.D(\buffer_9[17] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[17]_net_1 ));
    DFN1E1C0 \cur_scheme[33]  (.D(\buffer[34]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[33]));
    DFN1E1C0 \cur_flag[0]  (.D(\buffer[1]_net_1 ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(cur_flag_1_sqmuxa), .Q(
        demodulator_0_cur_flag[0]));
    DFN1E1C0 \cur_scheme[31]  (.D(\buffer[32]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[31]));
    NOR2A \buffer_RNO[37]  (.A(\buffer[36]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[37] ));
    DFN1E0C0 \buffer[44]  (.D(\buffer_9[44] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[44]_net_1 ));
    NOR2A \buffer_RNO[27]  (.A(\buffer[26]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[27] ));
    OR3 \latency_RNIQ2V32[1]  (.A(un1_buffer21_3_i_i_o2_1), .B(
        un1_buffer21_3_i_i_o2_0), .C(N_48), .Y(un1_buffer21_3_i_i_o2_5)
        );
    NOR2B un1_len_1_I_28 (.A(\DWACT_ADD_CI_0_g_array_1[0] ), .B(
        \len[2]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12[0] ));
    DFN1C0 \counter[5]  (.D(\counter_3[5] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[5]_net_1 ));
    NOR2B \len_RNO[2]  (.A(I_23), .B(un1_len_1_sqmuxa), .Y(\len_10[2] )
        );
    DFN1E1C0 \cur_flag[6]  (.D(\buffer[7]_net_1 ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(cur_flag_1_sqmuxa), .Q(
        demodulator_0_cur_flag[6]));
    NOR2B \waittime_RNIUNTF[2]  (.A(waittime_c1), .B(
        \waittime[2]_net_1 ), .Y(waittime_c2));
    NOR3B \buffer_RNI0JBT[50]  (.A(\buffer[49]_net_1 ), .B(
        \buffer[50]_net_1 ), .C(checksum_net_1), .Y(
        cur_scheme_0_sqmuxa_1));
    DFN1E1C0 \cur_scheme[36]  (.D(\buffer[37]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[36]));
    DFN1E0C0 \buffer[22]  (.D(\buffer_9[22] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[22]_net_1 ));
    DFN1E0C0 \buffer[34]  (.D(\buffer_9[34] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[34]_net_1 ));
    OR3B \latency_RNIJ4KO1[4]  (.A(\latency[3]_net_1 ), .B(
        \latency[4]_net_1 ), .C(N_40), .Y(N_42));
    XOR2 un3_counter_I_9 (.A(N_4), .B(\counter[3]_net_1 ), .Y(I_9));
    XA1C \latency_RNO[9]  (.A(\latency[9]_net_1 ), .B(N_55), .C(N_278), 
        .Y(latency_n9));
    OR2B \len_RNIEDAL81[3]  (.A(\len_RNI2H48I[3]_net_1 ), .B(
        un1_working_2), .Y(un1_len_1_sqmuxa));
    NOR2A \buffer_RNO[13]  (.A(\buffer[12]_net_1 ), .B(un1_working_2_0)
        , .Y(\buffer_9[13] ));
    DFN1E1C0 \ctg[0]  (.D(cur_flag_1_sqmuxa_i), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(ord_1_sqmuxa), .Q(demodulator_0_ctg[0]));
    NOR3B \buffer_RNIK8A3B[1]  (.A(ord34), .B(N_75_1), .C(ord10), .Y(
        len_3_sqmuxa_1));
    DFN1E0C0 \latency[1]  (.D(N_33), .CLK(ref_signal_c), .CLR(reset_c), 
        .E(N_8), .Q(\latency[1]_net_1 ));
    AND2 un1_len_1_I_35 (.A(\len[2]_net_1 ), .B(\len[3]_net_1 ), .Y(
        \DWACT_ADD_CI_0_pog_array_1[0] ));
    DFN1E0C0 \waittime[10]  (.D(waittime_n10), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(N_37), .Q(\waittime[10]_net_1 ));
    NOR2 \len_RNI2H48I[3]  (.A(un1_counter11_0), .B(len_3_sqmuxa), .Y(
        \len_RNI2H48I[3]_net_1 ));
    NOR2B \waittime_RNIPVJA[2]  (.A(\waittime[5]_net_1 ), .B(
        \waittime[2]_net_1 ), .Y(buffer21_4));
    NOR2A \buffer_RNO[43]  (.A(\buffer[42]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[43] ));
    NOR3B \len_RNIO6I0H[3]  (.A(buffer_3_sqmuxa_2), .B(
        len_3_sqmuxa_1_0), .C(ord34), .Y(len_3_sqmuxa));
    XOR2 un1_len_1_I_17 (.A(\len[0]_net_1 ), .B(
        \len_RNI2H48I[3]_net_1 ), .Y(\DWACT_ADD_CI_0_partial_sum[0] ));
    DFN1E0C0 \buffer[7]  (.D(\buffer_9[7] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(un1_counter11_0_0), .Q(\buffer[7]_net_1 ));
    XA1 \waittime_RNO[7]  (.A(waittime_c6), .B(\waittime[7]_net_1 ), 
        .C(latency_1_sqmuxa_1), .Y(waittime_n7));
    OR2 \latency_RNIFSKM[2]  (.A(\latency[2]_net_1 ), .B(
        \latency[3]_net_1 ), .Y(un1_LOWERBOUND_0lto9_2));
    OR2B \latency_RNICPKM[2]  (.A(\latency[2]_net_1 ), .B(
        \latency[0]_net_1 ), .Y(N_39));
    DFN1E1C0 \cur_scheme[42]  (.D(\buffer[43]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[42]));
    DFN1E0C0 \buffer[6]  (.D(\buffer_9[6] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(un1_counter11_0_0), .Q(\buffer[6]_net_1 ));
    XOR2 un3_counter_I_12 (.A(N_3), .B(\counter[4]_net_1 ), .Y(I_12));
    AX1A \latency_RNO_0[4]  (.A(N_40), .B(\latency[3]_net_1 ), .C(
        \latency[4]_net_1 ), .Y(latency_n4_i_0));
    DFN1E0C0 \buffer[19]  (.D(\buffer_9[19] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[19]_net_1 ));
    NOR2A \latency_RNIRHI7D[9]  (.A(un1_insig_i_0), .B(N_13), .Y(
        len_3_sqmuxa_1_0));
    NOR2 \latency_RNO[1]  (.A(latency_n1_i_0), .B(N_278), .Y(N_33));
    XOR2 ord_11_I_8 (.A(demodulator_0_ord[0]), .B(ord_1_sqmuxa), .Y(
        \DWACT_ADD_CI_0_partial_sum_0[0] ));
    DFN1E1C0 \cur_scheme[2]  (.D(\buffer[3]_net_1 ), .CLK(ref_signal_c)
        , .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[2]));
    DFN1E1C0 \cur_scheme[44]  (.D(\buffer[45]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[44]));
    OR2B \buffer_RNIOP0D1[1]  (.A(ord10), .B(ord34), .Y(ctg_0_sqmuxa));
    AO1A checksum_RNO (.A(N_58_i), .B(N_75_1), .C(checksum_4_iv_0_0), 
        .Y(checksum_4));
    NOR2A \buffer_RNO[16]  (.A(\buffer[15]_net_1 ), .B(un1_working_2_0)
        , .Y(\buffer_9[16] ));
    DFN1E1C0 \cur_scheme[1]  (.D(\buffer[2]_net_1 ), .CLK(ref_signal_c)
        , .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[1]));
    DFN1E1C0 \cur_flag[2]  (.D(\buffer[3]_net_1 ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(cur_flag_1_sqmuxa), .Q(
        demodulator_0_cur_flag[2]));
    NOR2B \waittime_RNIKR551[6]  (.A(waittime_c5), .B(
        \waittime[6]_net_1 ), .Y(waittime_c6));
    NOR2 \len_RNIHR87_0[5]  (.A(\len[5]_net_1 ), .B(\len[4]_net_1 ), 
        .Y(N_18));
    NOR2A \buffer_RNO[7]  (.A(\buffer[6]_net_1 ), .B(un1_working_2_0), 
        .Y(\buffer_9[7] ));
    XA1 \waittime_RNO[2]  (.A(waittime_c1), .B(\waittime[2]_net_1 ), 
        .C(latency_1_sqmuxa_1), .Y(waittime_n2));
    DFN1E1C0 \cur_scheme[15]  (.D(\buffer[16]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[15]));
    NOR2A \buffer_RNO[12]  (.A(\buffer[11]_net_1 ), .B(un1_working_2_0)
        , .Y(\buffer_9[12] ));
    DFN1E0C0 \buffer[47]  (.D(\buffer_9[47] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[47]_net_1 ));
    NOR3C \counter_RNID65O[1]  (.A(counter10_1), .B(counter10_0), .C(
        counter10_2), .Y(counter10));
    AO1 checksum_RNO_1 (.A(checksum_4_iv_0_a4_1_0), .B(buffer22), .C(
        N_76), .Y(checksum_4_iv_0_0));
    XOR2 un3_counter_I_7 (.A(N_5), .B(\counter[2]_net_1 ), .Y(I_7));
    OR2 \latency_RNIIDAD1[6]  (.A(un1_LOWERBOUND_0lto9_4), .B(
        un1_LOWERBOUND_0lto9_5), .Y(un1_LOWERBOUND_0lt9_1));
    XA1 \waittime_RNO[6]  (.A(waittime_c5), .B(\waittime[6]_net_1 ), 
        .C(latency_1_sqmuxa_1), .Y(waittime_n6));
    XOR2 un1_len_1_I_24 (.A(\len[1]_net_1 ), .B(
        \DWACT_ADD_CI_0_TMP[0] ), .Y(I_24));
    AO1 \counter_RNIRAAIH[1]  (.A(buffer_3_sqmuxa_2), .B(
        len_3_sqmuxa_1_0), .C(un1_counter11_0), .Y(un1_counter11_0_0));
    NOR2A \buffer_RNO[46]  (.A(\buffer[45]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[46] ));
    OR2 \latency_RNIERKM[1]  (.A(\latency[3]_net_1 ), .B(
        \latency[1]_net_1 ), .Y(un1_buffer21_3_i_i_o2_0));
    DFN1E1C0 \ctg[1]  (.D(ctg_0_sqmuxa), .CLK(ref_signal_c), .CLR(
        reset_c), .E(ord_1_sqmuxa), .Q(demodulator_0_ctg[1]));
    DFN1E0C0 \buffer[37]  (.D(\buffer_9[37] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[37]_net_1 ));
    NOR2A \buffer_RNO[42]  (.A(\buffer[41]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[42] ));
    DFN1E0C0 \waittime[0]  (.D(N_577), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_37), .Q(\waittime[0]_net_1 ));
    DFN1E0C0 \buffer[21]  (.D(\buffer_9[21] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[21]_net_1 ));
    DFN1E1C0 \cur_scheme[10]  (.D(\buffer[11]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[10]));
    DFN1E1C0 \cur_scheme[0]  (.D(\buffer[1]_net_1 ), .CLK(ref_signal_c)
        , .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[0]));
    NOR2A \buffer_RNO[15]  (.A(\buffer[14]_net_1 ), .B(un1_working_2_0)
        , .Y(\buffer_9[15] ));
    NOR3C \buffer_RNIFHTIF[50]  (.A(cur_scheme_0_sqmuxa), .B(counter10)
        , .C(len_3_sqmuxa_1_0), .Y(cur_scheme_1_sqmuxa));
    NOR3A \buffer_RNI8F5Q[9]  (.A(\buffer[10]_net_1 ), .B(
        \buffer[9]_net_1 ), .C(checksum_net_1), .Y(cur_flag_0_sqmuxa_1)
        );
    DFN1E0C0 \buffer[23]  (.D(\buffer_9[23] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[23]_net_1 ));
    NOR2B \waittime_RNI15A42[4]  (.A(buffer21_8), .B(buffer21_7), .Y(
        buffer21));
    DFN1E0C0 \buffer[12]  (.D(\buffer_9[12] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_0_0), .Q(\buffer[12]_net_1 ));
    DFN1E1C0 \cur_scheme[17]  (.D(\buffer[18]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[17]));
    NOR2A \counter_RNO[4]  (.A(I_12), .B(counter10), .Y(\counter_3[4] )
        );
    DFN1C0 \len[5]  (.D(\len_10[5] ), .CLK(ref_signal_c), .CLR(reset_c)
        , .Q(\len[5]_net_1 ));
    OR2 \latency_RNIN4LM[6]  (.A(\latency[7]_net_1 ), .B(
        \latency[6]_net_1 ), .Y(un1_LOWERBOUND_0lto9_4));
    NOR2A \buffer_RNO[45]  (.A(\buffer[44]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[45] ));
    NOR2B \waittime_RNI5PRV[5]  (.A(waittime_c4), .B(
        \waittime[5]_net_1 ), .Y(waittime_c5));
    XA1 \waittime_RNO[3]  (.A(waittime_c2), .B(\waittime[3]_net_1 ), 
        .C(latency_1_sqmuxa_1), .Y(waittime_n3));
    NOR3B \latency_RNIM0UFI[9]  (.A(un1_cur_scheme_0_sqmuxa), .B(
        ord_1_sqmuxa_0), .C(N_13), .Y(ord_1_sqmuxa));
    DFN1E0C0 \latency[0]  (.D(N_73), .CLK(ref_signal_c), .CLR(reset_c), 
        .E(N_8), .Q(\latency[0]_net_1 ));
    DFN1E0C0 \waittime[3]  (.D(waittime_n3), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_37), .Q(\waittime[3]_net_1 ));
    NOR2 \latency_RNO[5]  (.A(latency_n5_i_0), .B(N_278), .Y(N_25));
    NOR2A \buffer_RNO[38]  (.A(\buffer[37]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[38] ));
    DFN1E1C0 \cur_flag[4]  (.D(\buffer[5]_net_1 ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(cur_flag_1_sqmuxa), .Q(
        demodulator_0_cur_flag[4]));
    DFN1E0C0 \buffer[25]  (.D(\buffer_9[25] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[25]_net_1 ));
    XNOR2 \latency_RNO_0[1]  (.A(\latency[0]_net_1 ), .B(
        \latency[1]_net_1 ), .Y(latency_n1_i_0));
    NOR2A \buffer_RNO[28]  (.A(\buffer[27]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[28] ));
    OR2 \waittime_RNIU8NJ2_0[4]  (.A(checksum_0_sqmuxa), .B(
        mac_0_working), .Y(N_278));
    NOR2 un1_insig_i_0_a2 (.A(insig_c), .B(mac_0_working), .Y(
        un1_insig_i_0));
    DFN1C0 \len[2]  (.D(\len_10[2] ), .CLK(ref_signal_c), .CLR(reset_c)
        , .Q(\len[2]_net_1 ));
    OR2A \latency_RNIDLU32[5]  (.A(\latency[5]_net_1 ), .B(N_42), .Y(
        N_43));
    DFN1E1C0 \cur_flag[5]  (.D(\buffer[6]_net_1 ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(cur_flag_1_sqmuxa), .Q(
        demodulator_0_cur_flag[5]));
    NOR3C \buffer_RNIFHTIF_0[50]  (.A(cur_scheme_0_sqmuxa), .B(
        counter10), .C(len_3_sqmuxa_1_0), .Y(cur_scheme_1_sqmuxa_0));
    DFN1C0 \ord[1]  (.D(\ord_11[1] ), .CLK(ref_signal_c), .CLR(reset_c)
        , .Q(demodulator_0_ord[1]));
    DFN1E0C0 \buffer[49]  (.D(\buffer_9[49] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[49]_net_1 ));
    NOR2B un3_counter_I_11 (.A(\counter[3]_net_1 ), .B(
        \DWACT_FINC_E[0] ), .Y(N_3));
    NOR2B \len_RNO[5]  (.A(I_26), .B(un1_len_1_sqmuxa), .Y(\len_10[5] )
        );
    XOR2 un1_len_1_I_22 (.A(\len[3]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12[0] ), .Y(I_22));
    DFN1E1C0 \cur_scheme[29]  (.D(\buffer[30]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[29]));
    DFN1E0C0 \waittime[6]  (.D(waittime_n6), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_37), .Q(\waittime[6]_net_1 ));
    XOR2 \latency_RNO_0[3]  (.A(\latency[3]_net_1 ), .B(N_40), .Y(
        latency_n3_i_0));
    NOR2A \buffer_RNO[31]  (.A(\buffer[30]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[31] ));
    XOR2 \latency_RNO_0[5]  (.A(\latency[5]_net_1 ), .B(N_42), .Y(
        latency_n5_i_0));
    DFN1E1C0 \cur_flag[1]  (.D(\buffer[2]_net_1 ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(cur_flag_1_sqmuxa), .Q(
        demodulator_0_cur_flag[1]));
    NOR2A \buffer_RNO[21]  (.A(\buffer[20]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[21] ));
    DFN1E0C0 \buffer[39]  (.D(\buffer_9[39] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[39]_net_1 ));
    NOR3B checksum_RNO_3 (.A(insig_c), .B(checksum_net_1), .C(
        mac_0_working), .Y(N_76));
    DFN1E1C0 \cur_scheme[13]  (.D(\buffer[14]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[13]));
    DFN1E1C0 \cur_scheme[11]  (.D(\buffer[12]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[11]));
    OR3 \latency_RNIQK9D1[0]  (.A(\latency[0]_net_1 ), .B(
        \latency[1]_net_1 ), .C(un1_LOWERBOUND_0lto9_2), .Y(
        un1_LOWERBOUND_0lt9_0));
    DFN1E1C0 \cur_scheme[9]  (.D(\buffer[10]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[9]));
    MX2 \len_RNO[0]  (.A(len_3_sqmuxa_1), .B(
        \DWACT_ADD_CI_0_partial_sum[0] ), .S(un1_len_1_sqmuxa), .Y(
        \len_10[0] ));
    OR3 \latency_RNIV29H3[0]  (.A(un1_LOWERBOUND_0lt9_0), .B(N_48), .C(
        un1_LOWERBOUND_0lt9_1), .Y(un1_LOWERBOUND_0lto9));
    NOR2A \buffer_RNO[14]  (.A(\buffer[13]_net_1 ), .B(un1_working_2_0)
        , .Y(\buffer_9[14] ));
    NOR2A \waittime_RNO[0]  (.A(latency_1_sqmuxa_1), .B(
        \waittime[0]_net_1 ), .Y(N_577));
    AO1C \latency_RNO_0[2]  (.A(\latency[2]_net_1 ), .B(N_56), .C(N_40)
        , .Y(latency_n2_i_0));
    DFN1C0 \len[3]  (.D(\len_10[3] ), .CLK(ref_signal_c), .CLR(reset_c)
        , .Q(\len[3]_net_1 ));
    NOR3A \latency_RNIT5V32[0]  (.A(N_56), .B(un1_LOWERBOUND_0lto9_5), 
        .C(un1_LOWERBOUND_0lto9_4), .Y(un1_LOWERBOUND_0_1_2));
    DFN1E0C0 \buffer[4]  (.D(\buffer_9[4] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(un1_counter11_0_0), .Q(\buffer[4]_net_1 ));
    AO1 \latency_RNIVAS69_0[0]  (.A(un1_LOWERBOUND_0_1_3), .B(
        un1_LOWERBOUND_0lto9), .C(buffer21), .Y(un1_buffer21_1));
    OR2A \latency_RNI879F2[6]  (.A(\latency[6]_net_1 ), .B(N_43), .Y(
        N_44));
    DFN1E1C0 \cur_scheme[16]  (.D(\buffer[17]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[16]));
    DFN1E1C0 \cur_scheme[22]  (.D(\buffer[23]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[22]));
    NOR2A \buffer_RNO[6]  (.A(\buffer[5]_net_1 ), .B(un1_working_2_0), 
        .Y(\buffer_9[6] ));
    OR3A \buffer_RNIE86G4[1]  (.A(ctg_0_sqmuxa), .B(
        cur_scheme_0_sqmuxa), .C(cur_flag_0_sqmuxa), .Y(
        un1_cur_scheme_0_sqmuxa));
    NOR3A \buffer_RNIHJ6N[1]  (.A(\buffer[1]_net_1 ), .B(
        \buffer[2]_net_1 ), .C(checksum_net_1), .Y(ord10));
    NOR2A \buffer_RNO[10]  (.A(\buffer[9]_net_1 ), .B(un1_working_2_0), 
        .Y(\buffer_9[10] ));
    NOR2B \buffer_RNI7P5J1[50]  (.A(cur_scheme_0_sqmuxa_1), .B(ord36), 
        .Y(cur_scheme_0_sqmuxa));
    DFN1E1C0 \cur_scheme[24]  (.D(\buffer[25]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[24]));
    NOR2A \buffer_RNO[44]  (.A(\buffer[43]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[44] ));
    DFN1E1C0 \cur_scheme[39]  (.D(\buffer[40]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[39]));
    NOR2B \len_RNIO7TA[3]  (.A(\len[3]_net_1 ), .B(N_18), .Y(
        ord35_0_a2_0));
    AO1 \counter_RNIRAAIH_1[1]  (.A(buffer_3_sqmuxa_2), .B(
        len_3_sqmuxa_1_0), .C(un1_counter11_0), .Y(un1_counter11));
    DFN1E0C0 \buffer[20]  (.D(\buffer_9[20] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[20]_net_1 ));
    XA1C \latency_RNO[6]  (.A(\latency[6]_net_1 ), .B(N_43), .C(N_278), 
        .Y(N_23));
    INV \ctg_RNO[0]  (.A(cur_flag_1_sqmuxa), .Y(cur_flag_1_sqmuxa_i));
    NOR2B un1_len_1_I_33 (.A(\DWACT_ADD_CI_0_g_array_1[0] ), .B(
        \DWACT_ADD_CI_0_pog_array_1[0] ), .Y(
        \DWACT_ADD_CI_0_g_array_2[0] ));
    XOR2 un1_len_1_I_21 (.A(\len[4]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_2[0] ), .Y(I_21));
    DFN1E1C0 \cur_scheme[28]  (.D(\buffer[29]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[28]));
    MX2 \len_RNO[1]  (.A(len_3_sqmuxa_1), .B(I_24), .S(
        un1_len_1_sqmuxa), .Y(\len_10[1] ));
    DFN1E0C0 \buffer[42]  (.D(\buffer_9[42] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11), .Q(\buffer[42]_net_1 ));
    DFN1E1C0 \cur_flag[3]  (.D(\buffer[4]_net_1 ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(cur_flag_1_sqmuxa), .Q(
        demodulator_0_cur_flag[3]));
    DFN1E0C0 \waittime[9]  (.D(waittime_n9), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_37), .Q(\waittime[9]_net_1 ));
    NOR2A \buffer_RNO[40]  (.A(\buffer[39]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[40] ));
    DFN1E0C0 \buffer[11]  (.D(\buffer_9[11] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_0_0), .Q(\buffer[11]_net_1 ));
    NOR2B \len_RNO[4]  (.A(I_21), .B(un1_len_1_sqmuxa), .Y(\len_10[4] )
        );
    DFN1E0C0 \latency[4]  (.D(N_27), .CLK(ref_signal_c), .CLR(reset_c), 
        .E(N_8), .Q(\latency[4]_net_1 ));
    DFN1E0C0 \buffer[2]  (.D(\buffer_9[2] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(un1_counter11_0_0), .Q(\buffer[2]_net_1 ));
    DFN1E1C0 \cur_scheme[45]  (.D(\buffer[46]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[45]));
    OR2A \latency_RNICS5DM_1[9]  (.A(un1_buffer22), .B(mac_0_working), 
        .Y(un1_working_2_0));
    NOR2A \buffer_RNO[33]  (.A(\buffer[32]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[33] ));
    DFN1E0C0 \buffer[0]  (.D(checksum_2_sqmuxa), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_0_0), .Q(\buffer[0]_net_1 ));
    NOR2B \len_RNI76QL_1[3]  (.A(ord35_0_a2_0), .B(N_16), .Y(ord35));
    DFN1E0C0 \buffer[13]  (.D(\buffer_9[13] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_0_0), .Q(\buffer[13]_net_1 ));
    NOR2A \waittime_RNIQ0KA[8]  (.A(\waittime[8]_net_1 ), .B(
        \waittime[0]_net_1 ), .Y(buffer21_1));
    NOR2A \buffer_RNO[23]  (.A(\buffer[22]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[23] ));
    XA1C \latency_RNO[7]  (.A(\latency[7]_net_1 ), .B(N_44), .C(N_278), 
        .Y(N_21));
    OR3 \latency_RNI50AD1[9]  (.A(\latency[9]_net_1 ), .B(
        \latency[6]_net_1 ), .C(N_39), .Y(un1_buffer21_3_i_i_o2_4));
    DFN1E0C0 \buffer[32]  (.D(\buffer_9[32] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[32]_net_1 ));
    XA1 \waittime_RNO[1]  (.A(\waittime[1]_net_1 ), .B(
        \waittime[0]_net_1 ), .C(latency_1_sqmuxa_1), .Y(waittime_n1));
    NOR2 \latency_RNO[0]  (.A(\latency[0]_net_1 ), .B(N_278), .Y(N_73));
    DFN1E0C0 \waittime[8]  (.D(waittime_n8), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_37), .Q(\waittime[8]_net_1 ));
    DFN1E1C0 \cur_scheme[32]  (.D(\buffer[33]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa_0), .Q(
        demodulator_0_cur_scheme[32]));
    OR3 \len_RNIIBG0O[3]  (.A(buffer22), .B(waittimelde_i_o2_1), .C(
        N_79), .Y(N_61));
    DFN1E0C0 \buffer[8]  (.D(\buffer_9[8] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(un1_counter11_0_0), .Q(\buffer[8]_net_1 ));
    NOR2B \waittime_RNO_0[10]  (.A(\waittime[9]_net_1 ), .B(
        waittime_c8), .Y(waittime_22_0));
    NOR3B \waittime_RNIO58L[4]  (.A(\waittime[4]_net_1 ), .B(
        buffer21_4), .C(\waittime[9]_net_1 ), .Y(buffer21_7));
    DFN1C0 \ord[0]  (.D(\DWACT_ADD_CI_0_partial_sum_0[0] ), .CLK(
        ref_signal_c), .CLR(reset_c), .Q(demodulator_0_ord[0]));
    XA1C \latency_RNO[8]  (.A(\latency[8]_net_1 ), .B(N_54), .C(N_278), 
        .Y(N_19));
    DFN1E1C0 \cur_scheme[34]  (.D(\buffer[35]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[34]));
    DFN1E0C0 \waittime[4]  (.D(waittime_n4), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_37), .Q(\waittime[4]_net_1 ));
    DFN1E1C0 \cur_scheme[40]  (.D(\buffer[41]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[40]));
    DFN1E0C0 \buffer[15]  (.D(\buffer_9[15] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_0_0), .Q(\buffer[15]_net_1 ));
    NOR2B \waittime_RNINNHQ[4]  (.A(waittime_c3), .B(
        \waittime[4]_net_1 ), .Y(waittime_c4));
    DFN1E0C0 \latency[2]  (.D(N_31), .CLK(ref_signal_c), .CLR(reset_c), 
        .E(N_8), .Q(\latency[2]_net_1 ));
    DFN1E0C0 \buffer[26]  (.D(\buffer_9[26] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[26]_net_1 ));
    DFN1C0 \len[1]  (.D(\len_10[1] ), .CLK(ref_signal_c), .CLR(reset_c)
        , .Q(\len[1]_net_1 ));
    DFN1E1C0 \cur_scheme[38]  (.D(\buffer[39]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[38]));
    NOR2A \latency_RNISE9M9[0]  (.A(un1_insig_i_0), .B(un1_buffer21_1), 
        .Y(N_75_1));
    NOR2B \waittime_RNIAN7L[3]  (.A(waittime_c2), .B(
        \waittime[3]_net_1 ), .Y(waittime_c3));
    DFN1E1C0 \cur_scheme[47]  (.D(\buffer[48]_net_1 ), .CLK(
        ref_signal_c), .CLR(reset_c), .E(cur_scheme_1_sqmuxa), .Q(
        demodulator_0_cur_scheme[47]));
    NOR2A \buffer_RNO[19]  (.A(\buffer[18]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[19] ));
    DFN1E0C0 \buffer[28]  (.D(\buffer_9[28] ), .CLK(ref_signal_c), 
        .CLR(reset_c), .E(un1_counter11_1_0), .Q(\buffer[28]_net_1 ));
    DFN1E0C0 \latency[5]  (.D(N_25), .CLK(ref_signal_c), .CLR(reset_c), 
        .E(N_8), .Q(\latency[5]_net_1 ));
    NOR2 \latency_RNO[2]  (.A(latency_n2_i_0), .B(N_278), .Y(N_31));
    NOR2A \buffer_RNO[36]  (.A(\buffer[35]_net_1 ), .B(un1_working_2), 
        .Y(\buffer_9[36] ));
    OR3 \len_RNILIE12[3]  (.A(ord36), .B(ord35), .C(ord34), .Y(
        waittimelde_i_o2_1));
    AO1B \counter_RNITQCCR[1]  (.A(N_61), .B(latency_1_sqmuxa_1), .C(
        counter10), .Y(N_37));
    NOR2A \buffer_RNO[26]  (.A(\buffer[25]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[26] ));
    NOR2 \counter_RNIFN18[2]  (.A(\counter[2]_net_1 ), .B(
        \counter[3]_net_1 ), .Y(counter10_1));
    XOR2 un1_len_1_I_26 (.A(\len[5]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12_1[0] ), .Y(I_26));
    OR2 \latency_RNIP6LM[7]  (.A(\latency[8]_net_1 ), .B(
        \latency[7]_net_1 ), .Y(un1_buffer21_3_i_i_o2_1));
    DFN1C0 \counter[0]  (.D(I_4), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[0]_net_1 ));
    NOR2A \buffer_RNO[32]  (.A(\buffer[31]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[32] ));
    NOR2B \counter_RNIJR18[5]  (.A(\counter[5]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(counter10_0));
    OR2 \latency_RNIJ0LM[4]  (.A(\latency[5]_net_1 ), .B(
        \latency[4]_net_1 ), .Y(N_48));
    NOR2A \buffer_RNO[22]  (.A(\buffer[21]_net_1 ), .B(un1_working_2_1)
        , .Y(\buffer_9[22] ));
    DFN1E0C0 \buffer[1]  (.D(\buffer_9[1] ), .CLK(ref_signal_c), .CLR(
        reset_c), .E(un1_counter11_0_0), .Q(\buffer[1]_net_1 ));
    NOR2 \latency_RNO[3]  (.A(latency_n3_i_0), .B(N_278), .Y(N_29));
    
endmodule


module data_source(
       data_source_0_output_data,
       reset_c,
       ref_signal_c,
       mac_0_datacmd,
       mac_0_head,
       mac_0_sending,
       output_signal_c
    );
output data_source_0_output_data;
input  reset_c;
input  ref_signal_c;
input  mac_0_datacmd;
input  mac_0_head;
input  mac_0_sending;
input  output_signal_c;

    wire N_364, \counter_RNI419N3[1]_net_1 , N_703, 
        \counter_RNI6RP44[1]_net_1 , counter_n15_i_0, N_355, 
        counter_n13_i_0, N_356, counter_n15_i_a3_0_0, 
        \counter[14]_net_1 , \counter[15]_net_1 , counter_n11_i_0, 
        N_357, output_data_2_sqmuxa_i_o3_5, counter19_3, 
        output_data_2_sqmuxa_i_o3_0, output_data_2_sqmuxa_i_o3_4, 
        \counter[5]_net_1 , \counter[4]_net_1 , 
        output_data_2_sqmuxa_i_o3_2, counter19_4, \counter[1]_net_1 , 
        \counter[0]_net_1 , counter19_4_0, counter19_3_0, counter19_1, 
        counter19_14_0_o3_1, \counter[8]_net_1 , \counter[9]_net_1 , 
        N_702, N_701, N_372, N_337, counter_c7, N_373, N_339, N_367, 
        N_341, N_368, \counter[10]_net_1 , N_345, N_370, 
        \counter[12]_net_1 , N_361, N_351, N_700, N_347, N_699, N_343, 
        N_697, counter_n7, counter_c6, \counter[7]_net_1 , counter_n6, 
        \counter[6]_net_1 , counter_c5, counter_n5, counter_c4, 
        counter_n4, counter_c3, counter_n3, \counter[3]_net_1 , 
        counter_c2, counter_n2, \counter[2]_net_1 , counter_c1, 
        output_data_7, \state[143]_net_1 , N_353, N_335, 
        \state[72]_net_1 , N_692, N_333, \state[80]_net_1 , N_690, 
        N_331, \state[88]_net_1 , N_688, N_329, \state[74]_net_1 , 
        N_686, N_327, \state[82]_net_1 , N_684, N_325, 
        \state[90]_net_1 , N_682, N_323, \state[76]_net_1 , N_680, 
        N_321, \state[84]_net_1 , N_678, N_319, \state[92]_net_1 , 
        N_676, N_317, \state[78]_net_1 , N_674, N_315, 
        \state[86]_net_1 , N_672, N_313, \state[94]_net_1 , N_670, 
        N_311, \state[96]_net_1 , N_668, N_309, \state[99]_net_1 , 
        N_666, N_307, \state[102]_net_1 , N_664, N_305, 
        \state[64]_net_1 , N_662, \state_8[72] , \state[71]_net_1 , 
        N_660, \state_8[80] , \state[79]_net_1 , N_658, \state_8[88] , 
        \state[87]_net_1 , N_656, \state_8[74] , \state[73]_net_1 , 
        N_654, \state_8[82] , \state[81]_net_1 , N_652, \state_8[90] , 
        \state[89]_net_1 , N_650, \state_8[76] , \state[75]_net_1 , 
        N_648, \state_8[84] , \state[83]_net_1 , N_646, \state_8[92] , 
        \state[91]_net_1 , N_644, \state_8[78] , \state[77]_net_1 , 
        N_642, \state_8[86] , \state[85]_net_1 , N_640, \state_8[94] , 
        \state[93]_net_1 , N_638, \state_8[96] , \state[95]_net_1 , 
        N_636, \state_8[98] , \state[97]_net_1 , N_634, \state_8[99] , 
        \state[98]_net_1 , N_632, \state_8[101] , \state[100]_net_1 , 
        N_630, \state_8[102] , \state[101]_net_1 , N_628, 
        \state_8[64] , \state[63]_net_1 , N_626, \state_8[66] , 
        \state[65]_net_1 , N_624, \state_8[67] , \state[66]_net_1 , 
        N_622, \state_8[68] , \state[67]_net_1 , N_620, \state_8[69] , 
        \state[68]_net_1 , N_618, \state_8[70] , \state[69]_net_1 , 
        N_616, \state_8[71] , \state[70]_net_1 , N_614, N_135, 
        \state[104]_net_1 , N_612, N_133, \state[112]_net_1 , N_610, 
        N_131, \state[120]_net_1 , N_608, N_129, \state[128]_net_1 , 
        N_606, N_127, \state[136]_net_1 , N_604, N_125, 
        \state[107]_net_1 , N_602, N_123, \state[115]_net_1 , N_600, 
        N_121, \state[123]_net_1 , N_598, N_119, \state[131]_net_1 , 
        N_596, N_117, \state[139]_net_1 , N_594, N_115, 
        \state[110]_net_1 , N_592, N_113, \state[118]_net_1 , N_590, 
        N_111, \state[126]_net_1 , N_588, N_109, \state[134]_net_1 , 
        N_586, N_107, \state[142]_net_1 , N_584, \state_8[104] , 
        \state[103]_net_1 , N_582, \state_8[112] , \state[111]_net_1 , 
        N_580, \state_8[120] , \state[119]_net_1 , N_578, 
        \state_8[128] , \state[127]_net_1 , N_576, \state_8[136] , 
        \state[135]_net_1 , N_574, \state_8[106] , \state[105]_net_1 , 
        N_572, \state_8[114] , \state[113]_net_1 , N_570, 
        \state_8[122] , \state[121]_net_1 , N_568, \state_8[130] , 
        \state[129]_net_1 , N_566, \state_8[138] , \state[137]_net_1 , 
        N_564, \state_8[107] , \state[106]_net_1 , N_562, 
        \state_8[115] , \state[114]_net_1 , N_560, \state_8[123] , 
        \state[122]_net_1 , N_558, \state_8[131] , \state[130]_net_1 , 
        N_556, \state_8[139] , \state[138]_net_1 , N_554, 
        \state_8[109] , \state[108]_net_1 , N_552, \state_8[125] , 
        \state[124]_net_1 , N_533, \state_8[133] , \state[132]_net_1 , 
        N_531, \state_8[141] , \state[140]_net_1 , N_529, 
        \state_8[110] , \state[109]_net_1 , N_527, \state_8[118] , 
        \state[117]_net_1 , N_525, \state_8[126] , \state[125]_net_1 , 
        N_523, \state_8[134] , \state[133]_net_1 , N_521, 
        \state_8[142] , \state[141]_net_1 , N_519, N_80, 
        \state[24]_net_1 , N_517, N_78, \state[32]_net_1 , N_515, N_76, 
        \state[40]_net_1 , N_513, N_74, \state[27]_net_1 , N_511, N_72, 
        \state[35]_net_1 , N_509, N_70, \state[43]_net_1 , N_507, N_68, 
        \state[30]_net_1 , N_505, N_66, \state[38]_net_1 , N_503, N_64, 
        \state[46]_net_1 , N_501, N_62, \state[48]_net_1 , N_499, N_60, 
        \state[56]_net_1 , N_497, \state_8[24] , \state[23]_net_1 , 
        N_495, \state_8[32] , \state[31]_net_1 , N_493, \state_8[40] , 
        \state[39]_net_1 , N_491, \state_8[34] , \state[33]_net_1 , 
        N_487, \state_8[42] , \state[41]_net_1 , N_485, \state_8[35] , 
        \state[34]_net_1 , N_546, \state_8[43] , \state[42]_net_1 , 
        N_544, \state_8[29] , \state[28]_net_1 , N_542, \state_8[37] , 
        \state[36]_net_1 , N_540, \state_8[45] , \state[44]_net_1 , 
        N_538, \state_8[30] , \state[29]_net_1 , N_536, \state_8[38] , 
        \state[37]_net_1 , N_453, \state_8[46] , \state[45]_net_1 , 
        N_451, \state_8[48] , \state[47]_net_1 , N_449, \state_8[56] , 
        \state[55]_net_1 , N_447, \state_8[50] , \state[49]_net_1 , 
        N_445, \state_8[58] , \state[57]_net_1 , N_443, \state_8[51] , 
        \state[50]_net_1 , N_441, \state_8[59] , \state[58]_net_1 , 
        N_439, \state_8[52] , \state[51]_net_1 , N_437, \state_8[60] , 
        \state[59]_net_1 , N_435, \state_8[53] , \state[52]_net_1 , 
        N_433, \state_8[61] , \state[60]_net_1 , N_431, \state_8[54] , 
        \state[53]_net_1 , N_429, \state_8[62] , \state[61]_net_1 , 
        N_427, \state_8[55] , \state[54]_net_1 , N_425, \state_8[63] , 
        \state[62]_net_1 , N_423, \state_8[23] , \state[22]_net_1 , 
        N_421, \state_8[22] , \state[21]_net_1 , N_419, \state_8[21] , 
        \state[20]_net_1 , N_417, \state_8[20] , \state[19]_net_1 , 
        N_415, \state_8[19] , \state[18]_net_1 , N_413, \state_8[18] , 
        \state[17]_net_1 , N_411, \state_8[9] , \state[8]_net_1 , 
        N_393, \state_8[8] , \state[7]_net_1 , N_391, \state_8[7] , 
        \state[6]_net_1 , N_389, \state_8[6] , \state[5]_net_1 , N_387, 
        \state_8[5] , \state[4]_net_1 , N_385, \state_8[1] , 
        \state[0]_net_1 , N_377, \state_8[0] , N_375, 
        \state[116]_net_1 , \state[25]_net_1 , \state[9]_net_1 , 
        \state[1]_net_1 , counter_n1, counter_n0, N_379, 
        \state[2]_net_1 , N_381, \state[3]_net_1 , N_383, N_395, 
        \state[10]_net_1 , N_397, \state[11]_net_1 , N_399, 
        \state[12]_net_1 , N_401, \state[13]_net_1 , N_403, 
        \state[14]_net_1 , N_405, \state[15]_net_1 , N_407, 
        \state[16]_net_1 , N_409, N_483, N_489, \state[26]_net_1 , 
        N_550, \counter[11]_net_1 , \counter[13]_net_1 , \state_8[2] , 
        \state_8[3] , \state_8[4] , \state_8[10] , \state_8[11] , 
        \state_8[12] , \state_8[13] , \state_8[14] , \state_8[15] , 
        \state_8[16] , \state_8[17] , \state_8[27] , \state_8[26] , 
        \state_8[117] , N_349, N_369, N_371, GND, VCC;
    
    NOR3B \state_RNO_0[31]  (.A(output_signal_c), .B(N_364), .C(
        \state[31]_net_1 ), .Y(N_505));
    AO1 \state_RNO[27]  (.A(\state[26]_net_1 ), .B(N_703), .C(N_483), 
        .Y(\state_8[27] ));
    DFN1C0 \state[40]  (.D(\state_8[40] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[40]_net_1 ));
    DFN1P0 \state[111]  (.D(N_115), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[111]_net_1 ));
    NOR3B \state_RNO_0[91]  (.A(output_signal_c), .B(N_364), .C(
        \state[91]_net_1 ), .Y(N_682));
    NOR3B \state_RNO_0[44]  (.A(output_signal_c), .B(N_364), .C(
        \state[44]_net_1 ), .Y(N_507));
    NOR3C \state_RNO_0[29]  (.A(output_signal_c), .B(N_364), .C(
        \state[29]_net_1 ), .Y(N_542));
    DFN1C0 \state[0]  (.D(\state_8[0] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[0]_net_1 ));
    AO1 \state_RNO[136]  (.A(\state[135]_net_1 ), .B(N_703), .C(N_574), 
        .Y(\state_8[136] ));
    NOR3B \state_RNO_0[143]  (.A(output_signal_c), .B(N_364), .C(
        \state[143]_net_1 ), .Y(N_584));
    NOR3B \state_RNO_0[57]  (.A(output_signal_c), .B(N_364), .C(
        \state[57]_net_1 ), .Y(N_497));
    NOR3C \state_RNO_0[10]  (.A(output_signal_c), .B(N_364), .C(
        \state[10]_net_1 ), .Y(N_395));
    DFN1C0 \state[23]  (.D(\state_8[23] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[23]_net_1 ));
    NOR3C \state_RNO_0[37]  (.A(output_signal_c), .B(N_364), .C(
        \state[37]_net_1 ), .Y(N_540));
    NOR3C \state_RNO_0[20]  (.A(output_signal_c), .B(N_364), .C(
        \state[20]_net_1 ), .Y(N_415));
    NOR3B \state_RNO_0[97]  (.A(output_signal_c), .B(N_364), .C(
        \state[97]_net_1 ), .Y(N_668));
    DFN1C0 \state[114]  (.D(\state_8[114] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[114]_net_1 ));
    AO1 \state_RNO[22]  (.A(\state[21]_net_1 ), .B(N_703), .C(N_419), 
        .Y(\state_8[22] ));
    NOR3C \state_RNO_0[110]  (.A(output_signal_c), .B(N_364), .C(
        \state[110]_net_1 ), .Y(N_527));
    AO1 \state_RNO[43]  (.A(\state[42]_net_1 ), .B(N_703), .C(N_544), 
        .Y(\state_8[43] ));
    OR2 \counter_RNIVPDJ[1]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(output_data_2_sqmuxa_i_o3_0));
    AO1 \state_RNO[10]  (.A(\state[9]_net_1 ), .B(N_703), .C(N_395), 
        .Y(\state_8[10] ));
    DFN1C0 \state[29]  (.D(\state_8[29] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[29]_net_1 ));
    NOR3C \state_RNO_0[2]  (.A(output_signal_c), .B(N_364), .C(
        \state[2]_net_1 ), .Y(N_379));
    DFN1C0 \state[118]  (.D(\state_8[118] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[118]_net_1 ));
    NOR3C \state_RNO_0[52]  (.A(output_signal_c), .B(N_364), .C(
        \state[52]_net_1 ), .Y(N_437));
    AO1 \state_RNO[134]  (.A(\state[133]_net_1 ), .B(N_703), .C(N_521), 
        .Y(\state_8[134] ));
    DFN1C0 \state[55]  (.D(\state_8[55] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[55]_net_1 ));
    NOR2B \counter_RNI2OR61[3]  (.A(counter_c2), .B(\counter[3]_net_1 )
        , .Y(counter_c3));
    OA1C \state_RNO[95]  (.A(N_703), .B(\state[94]_net_1 ), .C(N_670), 
        .Y(N_313));
    NOR3C \state_RNO_0[32]  (.A(output_signal_c), .B(N_364), .C(
        \state[32]_net_1 ), .Y(N_493));
    AO1 \state_RNO[30]  (.A(\state[29]_net_1 ), .B(N_703), .C(N_536), 
        .Y(\state_8[30] ));
    NOR3A \counter_RNO[11]  (.A(N_370), .B(N_697), .C(counter_n11_i_0), 
        .Y(N_343));
    NOR3C \state_RNO_0[92]  (.A(output_signal_c), .B(N_364), .C(
        \state[92]_net_1 ), .Y(N_644));
    DFN1C0 \state[10]  (.D(\state_8[10] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[10]_net_1 ));
    AO1 \state_RNO[17]  (.A(\state[16]_net_1 ), .B(N_703), .C(N_409), 
        .Y(\state_8[17] ));
    DFN1P0 \state[81]  (.D(N_333), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[81]_net_1 ));
    NOR3C \state_RNO_0[136]  (.A(output_signal_c), .B(N_364), .C(
        \state[136]_net_1 ), .Y(N_574));
    AO1 \state_RNO[69]  (.A(\state[68]_net_1 ), .B(N_703), .C(N_618), 
        .Y(\state_8[69] ));
    DFN1P0 \state[57]  (.D(N_60), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[57]_net_1 ));
    DFN1C0 \counter[11]  (.D(N_343), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[11]_net_1 ));
    NOR3C \state_RNO_0[55]  (.A(output_signal_c), .B(N_364), .C(
        \state[55]_net_1 ), .Y(N_425));
    NOR3B \state_RNO_0[111]  (.A(output_signal_c), .B(N_364), .C(
        \state[111]_net_1 ), .Y(N_592));
    DFN1C0 \state[88]  (.D(\state_8[88] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[88]_net_1 ));
    DFN1C0 \state[6]  (.D(\state_8[6] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[6]_net_1 ));
    NOR3C \state_RNO_0[35]  (.A(output_signal_c), .B(N_364), .C(
        \state[35]_net_1 ), .Y(N_546));
    AO1 \state_RNO[37]  (.A(\state[36]_net_1 ), .B(N_703), .C(N_540), 
        .Y(\state_8[37] ));
    DFN1C0 \state[64]  (.D(\state_8[64] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[64]_net_1 ));
    NOR2B \counter_RNIGO4T[2]  (.A(counter_c1), .B(\counter[2]_net_1 ), 
        .Y(counter_c2));
    CLKINT \counter_RNI6RP44_0[1]  (.A(\counter_RNI6RP44[1]_net_1 ), 
        .Y(N_703));
    NOR3B \state_RNO_0[95]  (.A(output_signal_c), .B(N_364), .C(
        \state[95]_net_1 ), .Y(N_670));
    OA1C \state_RNO[113]  (.A(N_703), .B(\state[112]_net_1 ), .C(N_610)
        , .Y(N_133));
    NOR3 \counter_RNO[15]  (.A(N_700), .B(counter_n15_i_0), .C(N_701), 
        .Y(N_351));
    NOR3C \state_RNO_0[48]  (.A(output_signal_c), .B(N_364), .C(
        \state[48]_net_1 ), .Y(N_449));
    DFN1P0 \state[132]  (.D(N_119), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[132]_net_1 ));
    CLKINT \counter_RNI419N3_0[1]  (.A(\counter_RNI419N3[1]_net_1 ), 
        .Y(N_364));
    AO1 \state_RNO[123]  (.A(\state[122]_net_1 ), .B(N_703), .C(N_558), 
        .Y(\state_8[123] ));
    AO1 \state_RNO[12]  (.A(\state[11]_net_1 ), .B(N_703), .C(N_399), 
        .Y(\state_8[12] ));
    NOR3B \state_RNO_0[49]  (.A(output_signal_c), .B(N_364), .C(
        \state[49]_net_1 ), .Y(N_499));
    NOR3C \state_RNO_0[118]  (.A(output_signal_c), .B(N_364), .C(
        \state[118]_net_1 ), .Y(N_525));
    DFN1C0 \state[96]  (.D(\state_8[96] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[96]_net_1 ));
    AO1 \state_RNO[76]  (.A(\state[75]_net_1 ), .B(N_703), .C(N_648), 
        .Y(\state_8[76] ));
    OA1C \state_RNO[103]  (.A(N_703), .B(\state[102]_net_1 ), .C(N_664)
        , .Y(N_307));
    AO1 \state_RNO[56]  (.A(\state[55]_net_1 ), .B(N_703), .C(N_447), 
        .Y(\state_8[56] ));
    DFN1C0 \state[133]  (.D(\state_8[133] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[133]_net_1 ));
    NOR3C \state_RNO_0[40]  (.A(output_signal_c), .B(N_364), .C(
        \state[40]_net_1 ), .Y(N_491));
    OA1C \state_RNO[49]  (.A(N_703), .B(\state[48]_net_1 ), .C(N_499), 
        .Y(N_62));
    AO1 \state_RNO[32]  (.A(\state[31]_net_1 ), .B(N_703), .C(N_493), 
        .Y(\state_8[32] ));
    XA1B \counter_RNO[7]  (.A(counter_c6), .B(\counter[7]_net_1 ), .C(
        N_373), .Y(counter_n7));
    NOR3B \state_RNO_0[132]  (.A(output_signal_c), .B(N_364), .C(
        \state[132]_net_1 ), .Y(N_596));
    AO1 \state_RNO[80]  (.A(\state[79]_net_1 ), .B(N_703), .C(N_658), 
        .Y(\state_8[80] ));
    DFN1C0 \counter[6]  (.D(counter_n6), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[6]_net_1 ));
    DFN1C0 \state[102]  (.D(\state_8[102] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[102]_net_1 ));
    DFN1P0 \state[31]  (.D(N_68), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[31]_net_1 ));
    NOR2 \counter_RNIB6EJ[6]  (.A(\counter[6]_net_1 ), .B(
        \counter[7]_net_1 ), .Y(counter19_4));
    NOR3C \state_RNO_0[54]  (.A(output_signal_c), .B(N_364), .C(
        \state[54]_net_1 ), .Y(N_429));
    OR2 \counter_RNI5961[12]  (.A(\counter[13]_net_1 ), .B(
        \counter[12]_net_1 ), .Y(N_356));
    NOR3C \state_RNO_0[66]  (.A(output_signal_c), .B(N_364), .C(
        \state[66]_net_1 ), .Y(N_624));
    DFN1P0 \state[93]  (.D(N_319), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[93]_net_1 ));
    DFN1C0 \state[50]  (.D(\state_8[50] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[50]_net_1 ));
    DFN1C0 \state[38]  (.D(\state_8[38] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[38]_net_1 ));
    NOR3C \state_RNO_0[34]  (.A(output_signal_c), .B(N_364), .C(
        \state[34]_net_1 ), .Y(N_487));
    DFN1P0 \state[44]  (.D(N_70), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[44]_net_1 ));
    NOR3C \state_RNO_0[142]  (.A(output_signal_c), .B(N_364), .C(
        \state[142]_net_1 ), .Y(N_519));
    NOR3C \state_RNO_0[94]  (.A(output_signal_c), .B(N_364), .C(
        \state[94]_net_1 ), .Y(N_638));
    OAI1 output_data_RNO_0 (.A(N_361), .B(output_data_2_sqmuxa_i_o3_5), 
        .C(output_signal_c), .Y(N_353));
    DFN1C0 \counter[3]  (.D(counter_n3), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[3]_net_1 ));
    DFN1C0 \counter[2]  (.D(counter_n2), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[2]_net_1 ));
    AO1 \state_RNO[98]  (.A(\state[97]_net_1 ), .B(N_703), .C(N_634), 
        .Y(\state_8[98] ));
    DFN1P0 \state[103]  (.D(N_307), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[103]_net_1 ));
    XA1B \counter_RNO[8]  (.A(\counter[8]_net_1 ), .B(counter_c7), .C(
        N_373), .Y(N_337));
    AO1C \counter_RNIK0AI3[4]  (.A(N_361), .B(counter19_4_0), .C(
        output_signal_c), .Y(N_373));
    OA1C \state_RNO[87]  (.A(N_703), .B(\state[86]_net_1 ), .C(N_672), 
        .Y(N_315));
    NOR3A \counter_RNO[13]  (.A(N_372), .B(N_699), .C(counter_n13_i_0), 
        .Y(N_347));
    NOR2A \counter_RNO_0[11]  (.A(N_368), .B(\counter[11]_net_1 ), .Y(
        N_697));
    NOR2A \counter_RNI6RP44[1]  (.A(output_signal_c), .B(N_364), .Y(
        \counter_RNI6RP44[1]_net_1 ));
    NOR3C \state_RNO_0[115]  (.A(output_signal_c), .B(N_364), .C(
        \state[115]_net_1 ), .Y(N_560));
    DFN1C0 \state[99]  (.D(\state_8[99] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[99]_net_1 ));
    DFN1P0 \state[85]  (.D(N_321), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[85]_net_1 ));
    DFN1C0 \state[4]  (.D(\state_8[4] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[4]_net_1 ));
    NOR3C \state_RNO_0[71]  (.A(output_signal_c), .B(N_364), .C(
        \state[71]_net_1 ), .Y(N_614));
    NOR3B output_data_RNO_1 (.A(mac_0_head), .B(output_signal_c), .C(
        mac_0_datacmd), .Y(N_702));
    DFN1P0 \state[87]  (.D(N_315), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[87]_net_1 ));
    AO1 \state_RNO[82]  (.A(\state[81]_net_1 ), .B(N_703), .C(N_652), 
        .Y(\state_8[82] ));
    XA1C \counter_RNO[12]  (.A(N_370), .B(\counter[12]_net_1 ), .C(
        N_373), .Y(N_345));
    AO1 \state_RNO[115]  (.A(\state[114]_net_1 ), .B(N_703), .C(N_560), 
        .Y(\state_8[115] ));
    DFN1C0 \state[122]  (.D(\state_8[122] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[122]_net_1 ));
    AO1 \state_RNO[64]  (.A(\state[63]_net_1 ), .B(N_703), .C(N_626), 
        .Y(\state_8[64] ));
    DFN1C0 \state[7]  (.D(\state_8[7] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[7]_net_1 ));
    AO1 \state_RNO[26]  (.A(\state[25]_net_1 ), .B(N_703), .C(N_489), 
        .Y(\state_8[26] ));
    NOR3B \state_RNO_0[77]  (.A(output_signal_c), .B(N_364), .C(
        \state[77]_net_1 ), .Y(N_680));
    AO1 \state_RNO[125]  (.A(\state[124]_net_1 ), .B(N_703), .C(N_533), 
        .Y(\state_8[125] ));
    XA1B \counter_RNO[1]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .C(N_373), .Y(counter_n1));
    OR2 \counter_RNI9D61[14]  (.A(\counter[14]_net_1 ), .B(
        \counter[15]_net_1 ), .Y(N_355));
    DFN1C0 \state[14]  (.D(\state_8[14] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[14]_net_1 ));
    DFN1C0 \counter[4]  (.D(counter_n4), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[4]_net_1 ));
    DFN1C0 \state[5]  (.D(\state_8[5] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[5]_net_1 ));
    DFN1C0 \state[123]  (.D(\state_8[123] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[123]_net_1 ));
    DFN1C0 \counter[10]  (.D(N_341), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[10]_net_1 ));
    NOR3C \state_RNO_0[63]  (.A(output_signal_c), .B(N_364), .C(
        \state[63]_net_1 ), .Y(N_423));
    OA1C \state_RNO[105]  (.A(N_703), .B(\state[104]_net_1 ), .C(N_612)
        , .Y(N_135));
    NOR3C \state_RNO_0[58]  (.A(output_signal_c), .B(N_364), .C(
        \state[58]_net_1 ), .Y(N_443));
    DFN1C0 \state[136]  (.D(\state_8[136] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[136]_net_1 ));
    DFN1C0 \state[62]  (.D(\state_8[62] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[62]_net_1 ));
    AO1 \state_RNO[142]  (.A(\state[141]_net_1 ), .B(N_703), .C(N_519), 
        .Y(\state_8[142] ));
    GND GND_i (.Y(GND));
    DFN1C0 \counter[13]  (.D(N_347), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[13]_net_1 ));
    NOR3C \state_RNO_0[59]  (.A(output_signal_c), .B(N_364), .C(
        \state[59]_net_1 ), .Y(N_439));
    NOR3C \state_RNO_0[38]  (.A(output_signal_c), .B(N_364), .C(
        \state[38]_net_1 ), .Y(N_453));
    DFN1C0 \state[35]  (.D(\state_8[35] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[35]_net_1 ));
    DFN1P0 \state[140]  (.D(N_117), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[140]_net_1 ));
    NOR3C \state_RNO_0[72]  (.A(output_signal_c), .B(N_364), .C(
        \state[72]_net_1 ), .Y(N_660));
    NOR3C \state_RNO_0[98]  (.A(output_signal_c), .B(N_364), .C(
        \state[98]_net_1 ), .Y(N_634));
    NOR3B \state_RNO_0[39]  (.A(output_signal_c), .B(N_364), .C(
        \state[39]_net_1 ), .Y(N_503));
    OA1C \state_RNO[44]  (.A(N_703), .B(\state[43]_net_1 ), .C(N_507), 
        .Y(N_70));
    NOR3C \state_RNO_0[99]  (.A(output_signal_c), .B(N_364), .C(
        \state[99]_net_1 ), .Y(N_632));
    NOR3C \state_RNO_0[50]  (.A(output_signal_c), .B(N_364), .C(
        \state[50]_net_1 ), .Y(N_445));
    DFN1C0 \counter[12]  (.D(N_345), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[12]_net_1 ));
    NOR3C \state_RNO_0[5]  (.A(output_signal_c), .B(N_364), .C(
        \state[5]_net_1 ), .Y(N_385));
    NOR3C \state_RNO_0[4]  (.A(output_signal_c), .B(N_364), .C(
        \state[4]_net_1 ), .Y(N_383));
    DFN1C0 \state[37]  (.D(\state_8[37] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[37]_net_1 ));
    OA1C \state_RNO[65]  (.A(N_703), .B(\state[64]_net_1 ), .C(N_662), 
        .Y(N_305));
    NOR3C \state_RNO_0[130]  (.A(output_signal_c), .B(N_364), .C(
        \state[130]_net_1 ), .Y(N_566));
    AO1 \state_RNO[71]  (.A(\state[70]_net_1 ), .B(N_703), .C(N_614), 
        .Y(\state_8[71] ));
    NOR3C \state_RNO_0[30]  (.A(output_signal_c), .B(N_364), .C(
        \state[30]_net_1 ), .Y(N_536));
    DFN1C0 \state[80]  (.D(\state_8[80] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[80]_net_1 ));
    DFN1C0 \state[106]  (.D(\state_8[106] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[106]_net_1 ));
    NOR3B \state_RNO_0[75]  (.A(output_signal_c), .B(N_364), .C(
        \state[75]_net_1 ), .Y(N_686));
    AO1 \state_RNO[51]  (.A(\state[50]_net_1 ), .B(N_703), .C(N_441), 
        .Y(\state_8[51] ));
    NOR3C \state_RNO_0[90]  (.A(output_signal_c), .B(N_364), .C(
        \state[90]_net_1 ), .Y(N_650));
    NOR3C \state_RNO_0[7]  (.A(output_signal_c), .B(N_364), .C(
        \state[7]_net_1 ), .Y(N_389));
    AO1 \state_RNO[16]  (.A(\state[15]_net_1 ), .B(N_703), .C(N_407), 
        .Y(\state_8[16] ));
    AO1 \state_RNO[118]  (.A(\state[117]_net_1 ), .B(N_703), .C(N_525), 
        .Y(\state_8[118] ));
    DFN1C0 \state[71]  (.D(\state_8[71] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[71]_net_1 ));
    AO1 \state_RNO[128]  (.A(\state[127]_net_1 ), .B(N_703), .C(N_576), 
        .Y(\state_8[128] ));
    OR2B \counter_RNI1Q101[6]  (.A(mac_0_sending), .B(counter19_4), .Y(
        output_data_2_sqmuxa_i_o3_2));
    NOR3B \state_RNO_0[140]  (.A(output_signal_c), .B(N_364), .C(
        \state[140]_net_1 ), .Y(N_594));
    DFN1C0 \state[78]  (.D(\state_8[78] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[78]_net_1 ));
    OA1C \state_RNO[140]  (.A(N_703), .B(\state[139]_net_1 ), .C(N_594)
        , .Y(N_117));
    DFN1C0 \state[42]  (.D(\state_8[42] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[42]_net_1 ));
    OA1C \state_RNO[36]  (.A(N_703), .B(\state[35]_net_1 ), .C(N_509), 
        .Y(N_72));
    DFN1C0 \state[54]  (.D(\state_8[54] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[54]_net_1 ));
    NOR3B \state_RNO_0[129]  (.A(output_signal_c), .B(N_364), .C(
        \state[129]_net_1 ), .Y(N_606));
    OA1C \state_RNO[108]  (.A(N_703), .B(\state[107]_net_1 ), .C(N_602)
        , .Y(N_125));
    OR2B \counter_RNO_1[11]  (.A(N_357), .B(output_signal_c), .Y(
        counter_n11_i_0));
    NOR3C \state_RNO_0[86]  (.A(output_signal_c), .B(N_364), .C(
        \state[86]_net_1 ), .Y(N_640));
    AO1 \state_RNO[90]  (.A(\state[89]_net_1 ), .B(N_703), .C(N_650), 
        .Y(\state_8[90] ));
    NOR3C \state_RNO_0[131]  (.A(output_signal_c), .B(N_364), .C(
        \state[131]_net_1 ), .Y(N_556));
    OR2A \counter_RNI3B613[9]  (.A(\counter[9]_net_1 ), .B(N_367), .Y(
        N_368));
    OA1C \state_RNO[73]  (.A(N_703), .B(\state[72]_net_1 ), .C(N_692), 
        .Y(N_335));
    AO1 \state_RNO[45]  (.A(\state[44]_net_1 ), .B(N_703), .C(N_538), 
        .Y(\state_8[45] ));
    NOR3C \state_RNO_0[109]  (.A(output_signal_c), .B(N_364), .C(
        \state[109]_net_1 ), .Y(N_552));
    AO1 \state_RNO[1]  (.A(\state[0]_net_1 ), .B(N_703), .C(N_377), .Y(
        \state_8[1] ));
    AO1 \state_RNO[53]  (.A(\state[52]_net_1 ), .B(N_703), .C(N_433), 
        .Y(\state_8[53] ));
    DFN1C0 \counter[15]  (.D(N_351), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[15]_net_1 ));
    OR3 \counter_RNIGFKK[8]  (.A(\counter[8]_net_1 ), .B(
        \counter[9]_net_1 ), .C(N_357), .Y(counter19_14_0_o3_1));
    NOR3C \state_RNO_0[141]  (.A(output_signal_c), .B(N_364), .C(
        \state[141]_net_1 ), .Y(N_529));
    NOR3C \state_RNO_0[74]  (.A(output_signal_c), .B(N_364), .C(
        \state[74]_net_1 ), .Y(N_654));
    DFN1C0 \state[126]  (.D(\state_8[126] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[126]_net_1 ));
    DFN1C0 \state[30]  (.D(\state_8[30] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[30]_net_1 ));
    DFN1C0 \state[21]  (.D(\state_8[21] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[21]_net_1 ));
    NOR3C \state_RNO_0[0]  (.A(output_signal_c), .B(N_364), .C(
        \state[0]_net_1 ), .Y(N_375));
    OA1C \state_RNO[97]  (.A(N_703), .B(\state[96]_net_1 ), .C(N_668), 
        .Y(N_311));
    NOR3C \state_RNO_0[138]  (.A(output_signal_c), .B(N_364), .C(
        \state[138]_net_1 ), .Y(N_564));
    AO1 output_data_RNO (.A(\state[143]_net_1 ), .B(N_703), .C(N_702), 
        .Y(output_data_7));
    DFN1P0 \state[28]  (.D(N_74), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[28]_net_1 ));
    OR2A \counter_RNI9PI33[13]  (.A(\counter[13]_net_1 ), .B(N_371), 
        .Y(N_372));
    DFN1C0 \state[66]  (.D(\state_8[66] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[66]_net_1 ));
    DFN1C0 \state[141]  (.D(\state_8[141] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[141]_net_1 ));
    AO1 \state_RNO[21]  (.A(\state[20]_net_1 ), .B(N_703), .C(N_417), 
        .Y(\state_8[21] ));
    DFN1C0 \state[12]  (.D(\state_8[12] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[12]_net_1 ));
    VCC VCC_i (.Y(VCC));
    XA1C \counter_RNO[14]  (.A(N_372), .B(\counter[14]_net_1 ), .C(
        N_373), .Y(N_349));
    AO1 \state_RNO[68]  (.A(\state[67]_net_1 ), .B(N_703), .C(N_620), 
        .Y(\state_8[68] ));
    AO1 \state_RNO[86]  (.A(\state[85]_net_1 ), .B(N_703), .C(N_640), 
        .Y(\state_8[86] ));
    DFN1C0 \counter[1]  (.D(counter_n1), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[1]_net_1 ));
    DFN1C0 \state[112]  (.D(\state_8[112] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[112]_net_1 ));
    AO1 \state_RNO[92]  (.A(\state[91]_net_1 ), .B(N_703), .C(N_644), 
        .Y(\state_8[92] ));
    AO1 \state_RNO[112]  (.A(\state[111]_net_1 ), .B(N_703), .C(N_580), 
        .Y(\state_8[112] ));
    XA1B \counter_RNO[5]  (.A(\counter[5]_net_1 ), .B(counter_c4), .C(
        N_373), .Y(counter_n5));
    AO1 \state_RNO[122]  (.A(\state[121]_net_1 ), .B(N_703), .C(N_568), 
        .Y(\state_8[122] ));
    DFN1P0 \state[75]  (.D(N_329), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[75]_net_1 ));
    DFN1C0 \state[63]  (.D(\state_8[63] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[63]_net_1 ));
    NOR3B \state_RNO_0[83]  (.A(output_signal_c), .B(N_364), .C(
        \state[83]_net_1 ), .Y(N_684));
    NOR2 \counter_RNI3UDJ[2]  (.A(\counter[2]_net_1 ), .B(
        \counter[3]_net_1 ), .Y(counter19_3));
    NOR3B \state_RNO_0[127]  (.A(output_signal_c), .B(N_364), .C(
        \state[127]_net_1 ), .Y(N_588));
    AO1 \state_RNO[4]  (.A(\state[3]_net_1 ), .B(N_703), .C(N_383), .Y(
        \state_8[4] ));
    XA1B \counter_RNO[3]  (.A(\counter[3]_net_1 ), .B(counter_c2), .C(
        N_373), .Y(counter_n3));
    NOR3C \state_RNO_0[16]  (.A(output_signal_c), .B(N_364), .C(
        \state[16]_net_1 ), .Y(N_407));
    DFN1P0 \state[113]  (.D(N_133), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[113]_net_1 ));
    NOR3B \state_RNO_0[124]  (.A(output_signal_c), .B(N_364), .C(
        \state[124]_net_1 ), .Y(N_598));
    NOR3C \state_RNO_0[123]  (.A(output_signal_c), .B(N_364), .C(
        \state[123]_net_1 ), .Y(N_558));
    AO1 \state_RNO[23]  (.A(\state[22]_net_1 ), .B(N_703), .C(N_421), 
        .Y(\state_8[23] ));
    AO1 \state_RNO[102]  (.A(\state[101]_net_1 ), .B(N_703), .C(N_628), 
        .Y(\state_8[102] ));
    DFN1P0 \state[77]  (.D(N_323), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[77]_net_1 ));
    NOR3C \state_RNO_0[26]  (.A(output_signal_c), .B(N_364), .C(
        \state[26]_net_1 ), .Y(N_489));
    NOR3B \state_RNO_0[135]  (.A(output_signal_c), .B(N_364), .C(
        \state[135]_net_1 ), .Y(N_586));
    OA1C \state_RNO[79]  (.A(N_703), .B(\state[78]_net_1 ), .C(N_674), 
        .Y(N_317));
    NOR3C \state_RNO_0[107]  (.A(output_signal_c), .B(N_364), .C(
        \state[107]_net_1 ), .Y(N_562));
    AO1 \state_RNO[59]  (.A(\state[58]_net_1 ), .B(N_703), .C(N_439), 
        .Y(\state_8[59] ));
    AO1 \state_RNO[141]  (.A(\state[140]_net_1 ), .B(N_703), .C(N_529), 
        .Y(\state_8[141] ));
    DFN1C0 \state[9]  (.D(\state_8[9] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[9]_net_1 ));
    DFN1C0 \state[46]  (.D(\state_8[46] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[46]_net_1 ));
    DFN1C0 \state[69]  (.D(\state_8[69] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[69]_net_1 ));
    AO1 \state_RNO[48]  (.A(\state[47]_net_1 ), .B(N_703), .C(N_449), 
        .Y(\state_8[48] ));
    AO1 \state_RNO[2]  (.A(\state[1]_net_1 ), .B(N_703), .C(N_379), .Y(
        \state_8[2] ));
    DFN1C0 \state[84]  (.D(\state_8[84] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[84]_net_1 ));
    NOR3C \state_RNO_0[104]  (.A(output_signal_c), .B(N_364), .C(
        \state[104]_net_1 ), .Y(N_582));
    NOR3B \state_RNO_0[103]  (.A(output_signal_c), .B(N_364), .C(
        \state[103]_net_1 ), .Y(N_664));
    DFN1C0 \counter[5]  (.D(counter_n5), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[5]_net_1 ));
    NOR3C \state_RNO_0[78]  (.A(output_signal_c), .B(N_364), .C(
        \state[78]_net_1 ), .Y(N_642));
    AO1 \state_RNO[11]  (.A(\state[10]_net_1 ), .B(N_703), .C(N_397), 
        .Y(\state_8[11] ));
    AO1 \state_RNO[110]  (.A(\state[109]_net_1 ), .B(N_703), .C(N_527), 
        .Y(\state_8[110] ));
    OR3 \counter_RNIU51N[8]  (.A(N_355), .B(N_356), .C(
        counter19_14_0_o3_1), .Y(N_361));
    NOR3B \state_RNO_0[79]  (.A(output_signal_c), .B(N_364), .C(
        \state[79]_net_1 ), .Y(N_674));
    AO1 \state_RNO[120]  (.A(\state[119]_net_1 ), .B(N_703), .C(N_578), 
        .Y(\state_8[120] ));
    DFN1C0 \state[52]  (.D(\state_8[52] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[52]_net_1 ));
    DFN1P0 \state[25]  (.D(N_80), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[25]_net_1 ));
    OA1C \state_RNO[31]  (.A(N_703), .B(\state[30]_net_1 ), .C(N_505), 
        .Y(N_68));
    AO1 \state_RNO[133]  (.A(\state[132]_net_1 ), .B(N_703), .C(N_531), 
        .Y(\state_8[133] ));
    DFN1C0 \state[43]  (.D(\state_8[43] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[43]_net_1 ));
    XA1C \counter_RNO[10]  (.A(N_368), .B(\counter[10]_net_1 ), .C(
        N_373), .Y(N_341));
    NOR3C \state_RNO_0[70]  (.A(output_signal_c), .B(N_364), .C(
        \state[70]_net_1 ), .Y(N_616));
    AO1 \state_RNO[6]  (.A(\state[5]_net_1 ), .B(N_703), .C(N_387), .Y(
        \state_8[6] ));
    OA1C \state_RNO[100]  (.A(N_703), .B(\state[99]_net_1 ), .C(N_666), 
        .Y(N_309));
    NOR3C \state_RNO_0[61]  (.A(output_signal_c), .B(N_364), .C(
        \state[61]_net_1 ), .Y(N_431));
    DFN1C0 \state[27]  (.D(\state_8[27] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[27]_net_1 ));
    DFN1P0 \state[91]  (.D(N_325), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[91]_net_1 ));
    DFN1P0 \state[49]  (.D(N_62), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[49]_net_1 ));
    AO1 \state_RNO[13]  (.A(\state[12]_net_1 ), .B(N_703), .C(N_401), 
        .Y(\state_8[13] ));
    DFN1C0 \state[16]  (.D(\state_8[16] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[16]_net_1 ));
    OR3A \counter_RNI419N3[1]  (.A(mac_0_datacmd), .B(N_361), .C(
        output_data_2_sqmuxa_i_o3_5), .Y(\counter_RNI419N3[1]_net_1 ));
    NOR3C \state_RNO_0[13]  (.A(output_signal_c), .B(N_364), .C(
        \state[13]_net_1 ), .Y(N_401));
    DFN1C0 \state[70]  (.D(\state_8[70] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[70]_net_1 ));
    DFN1P0 \state[135]  (.D(N_109), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[135]_net_1 ));
    DFN1C0 \state[98]  (.D(\state_8[98] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[98]_net_1 ));
    NOR3C \state_RNO_0[67]  (.A(output_signal_c), .B(N_364), .C(
        \state[67]_net_1 ), .Y(N_622));
    NOR3C \state_RNO_0[126]  (.A(output_signal_c), .B(N_364), .C(
        \state[126]_net_1 ), .Y(N_523));
    DFN1C0 \state[34]  (.D(\state_8[34] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[34]_net_1 ));
    NOR3C \state_RNO_0[23]  (.A(output_signal_c), .B(N_364), .C(
        \state[23]_net_1 ), .Y(N_421));
    AO1 \state_RNO[29]  (.A(\state[28]_net_1 ), .B(N_703), .C(N_542), 
        .Y(\state_8[29] ));
    OA1C \state_RNO[33]  (.A(N_703), .B(\state[32]_net_1 ), .C(N_515), 
        .Y(N_78));
    AO1 \state_RNO[7]  (.A(\state[6]_net_1 ), .B(N_703), .C(N_389), .Y(
        \state_8[7] ));
    OR2A \counter_RNI3DP13[10]  (.A(\counter[10]_net_1 ), .B(N_368), 
        .Y(N_369));
    NOR2A \counter_RNO_2[15]  (.A(counter_n15_i_a3_0_0), .B(N_372), .Y(
        N_701));
    NOR3C \state_RNO_0[106]  (.A(output_signal_c), .B(N_364), .C(
        \state[106]_net_1 ), .Y(N_572));
    DFN1P0 \state[116]  (.D(N_123), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[116]_net_1 ));
    NOR3C \state_RNO_0[46]  (.A(output_signal_c), .B(N_364), .C(
        \state[46]_net_1 ), .Y(N_451));
    DFN1C0 \state[13]  (.D(\state_8[13] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[13]_net_1 ));
    NOR3C \state_RNO_0[1]  (.A(output_signal_c), .B(N_364), .C(
        \state[1]_net_1 ), .Y(N_377));
    OR2 \counter_RNI1561[10]  (.A(\counter[11]_net_1 ), .B(
        \counter[10]_net_1 ), .Y(N_357));
    AO1 \state_RNO[60]  (.A(\state[59]_net_1 ), .B(N_703), .C(N_435), 
        .Y(\state_8[60] ));
    DFN1P0 \state[105]  (.D(N_135), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[105]_net_1 ));
    OA1C \state_RNO[81]  (.A(N_703), .B(\state[80]_net_1 ), .C(N_690), 
        .Y(N_333));
    NOR3C \state_RNO_0[62]  (.A(output_signal_c), .B(N_364), .C(
        \state[62]_net_1 ), .Y(N_427));
    NOR2B \counter_RNIVPDJ_0[1]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(counter_c1));
    XA1B \counter_RNO[6]  (.A(\counter[6]_net_1 ), .B(counter_c5), .C(
        N_373), .Y(counter_n6));
    NOR3C \state_RNO_0[9]  (.A(output_signal_c), .B(N_364), .C(
        \state[9]_net_1 ), .Y(N_393));
    NOR3C \counter_RNI6SR61[4]  (.A(\counter[4]_net_1 ), .B(
        \counter[0]_net_1 ), .C(counter19_1), .Y(counter19_3_0));
    DFN1C0 \state[8]  (.D(\state_8[8] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[8]_net_1 ));
    OR2B \counter_RNIB5FN2[8]  (.A(counter_c7), .B(\counter[8]_net_1 ), 
        .Y(N_367));
    AO1 \state_RNO[74]  (.A(\state[73]_net_1 ), .B(N_703), .C(N_654), 
        .Y(\state_8[74] ));
    DFN1C0 \state[20]  (.D(\state_8[20] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[20]_net_1 ));
    DFN1C0 \state[19]  (.D(\state_8[19] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[19]_net_1 ));
    AO1 \state_RNO[54]  (.A(\state[53]_net_1 ), .B(N_703), .C(N_429), 
        .Y(\state_8[54] ));
    NOR3C \state_RNO_0[122]  (.A(output_signal_c), .B(N_364), .C(
        \state[122]_net_1 ), .Y(N_568));
    AO1 \state_RNO[96]  (.A(\state[95]_net_1 ), .B(N_703), .C(N_636), 
        .Y(\state_8[96] ));
    AO1 \state_RNO[67]  (.A(\state[66]_net_1 ), .B(N_703), .C(N_622), 
        .Y(\state_8[67] ));
    NOR3B \state_RNO_0[65]  (.A(output_signal_c), .B(N_364), .C(
        \state[65]_net_1 ), .Y(N_662));
    OA1C \state_RNO[111]  (.A(N_703), .B(\state[110]_net_1 ), .C(N_592)
        , .Y(N_115));
    AO1 \state_RNO[117]  (.A(\state[116]_net_1 ), .B(N_703), .C(N_550), 
        .Y(\state_8[117] ));
    OA1C \state_RNO[135]  (.A(N_703), .B(\state[134]_net_1 ), .C(N_586)
        , .Y(N_109));
    OA1C \state_RNO[121]  (.A(N_703), .B(\state[120]_net_1 ), .C(N_608)
        , .Y(N_131));
    OA1C \state_RNO[127]  (.A(N_703), .B(\state[126]_net_1 ), .C(N_588)
        , .Y(N_111));
    OA1C \state_RNO[119]  (.A(N_703), .B(\state[118]_net_1 ), .C(N_590)
        , .Y(N_113));
    DFN1C0 \state[56]  (.D(\state_8[56] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[56]_net_1 ));
    NOR3C \state_RNO_0[102]  (.A(output_signal_c), .B(N_364), .C(
        \state[102]_net_1 ), .Y(N_628));
    DFN1C0 \state[82]  (.D(\state_8[82] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[82]_net_1 ));
    AO1 \state_RNO[19]  (.A(\state[18]_net_1 ), .B(N_703), .C(N_413), 
        .Y(\state_8[19] ));
    OA1C \state_RNO[129]  (.A(N_703), .B(\state[128]_net_1 ), .C(N_606)
        , .Y(N_129));
    DFN1P0 \state[137]  (.D(N_127), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[137]_net_1 ));
    OA1C \state_RNO[83]  (.A(N_703), .B(\state[82]_net_1 ), .C(N_684), 
        .Y(N_327));
    AO1 \state_RNO[40]  (.A(\state[39]_net_1 ), .B(N_703), .C(N_491), 
        .Y(\state_8[40] ));
    DFN1C0 \state[3]  (.D(\state_8[3] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[3]_net_1 ));
    AO1 \state_RNO[101]  (.A(\state[100]_net_1 ), .B(N_703), .C(N_630), 
        .Y(\state_8[101] ));
    DFN1P0 \state[95]  (.D(N_313), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[95]_net_1 ));
    DFN1C0 \counter[14]  (.D(N_349), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[14]_net_1 ));
    AO1 \state_RNO[107]  (.A(\state[106]_net_1 ), .B(N_703), .C(N_562), 
        .Y(\state_8[107] ));
    DFN1E1C0 output_data (.D(output_data_7), .CLK(ref_signal_c), .CLR(
        reset_c), .E(N_353), .Q(data_source_0_output_data));
    AO1 \state_RNO[62]  (.A(\state[61]_net_1 ), .B(N_703), .C(N_427), 
        .Y(\state_8[62] ));
    DFN1C0 \state[125]  (.D(\state_8[125] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[125]_net_1 ));
    OA1C \state_RNO[39]  (.A(N_703), .B(\state[38]_net_1 ), .C(N_503), 
        .Y(N_66));
    AO1 \state_RNO[109]  (.A(\state[108]_net_1 ), .B(N_703), .C(N_552), 
        .Y(\state_8[109] ));
    DFN1C0 \state[130]  (.D(\state_8[130] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[130]_net_1 ));
    NOR3C \state_RNO_0[43]  (.A(output_signal_c), .B(N_364), .C(
        \state[43]_net_1 ), .Y(N_544));
    DFN1C0 \state[53]  (.D(\state_8[53] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[53]_net_1 ));
    DFN1P0 \state[97]  (.D(N_311), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[97]_net_1 ));
    OA1C \state_RNO[75]  (.A(N_703), .B(\state[74]_net_1 ), .C(N_686), 
        .Y(N_329));
    OA1C \state_RNO[47]  (.A(N_703), .B(\state[46]_net_1 ), .C(N_501), 
        .Y(N_64));
    NOR2A \counter_RNO_0[13]  (.A(N_370), .B(\counter[13]_net_1 ), .Y(
        N_699));
    AO1 \state_RNO[55]  (.A(\state[54]_net_1 ), .B(N_703), .C(N_425), 
        .Y(\state_8[55] ));
    DFN1C0 \state[107]  (.D(\state_8[107] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[107]_net_1 ));
    NOR3C \state_RNO_0[64]  (.A(output_signal_c), .B(N_364), .C(
        \state[64]_net_1 ), .Y(N_626));
    DFN1C0 \state[139]  (.D(\state_8[139] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[139]_net_1 ));
    DFN1C0 \state[59]  (.D(\state_8[59] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[59]_net_1 ));
    NOR3B \state_RNO_0[81]  (.A(output_signal_c), .B(N_364), .C(
        \state[81]_net_1 ), .Y(N_690));
    AO1 \state_RNO[24]  (.A(\state[23]_net_1 ), .B(N_703), .C(N_495), 
        .Y(\state_8[24] ));
    OA1C \state_RNO[116]  (.A(N_703), .B(\state[115]_net_1 ), .C(N_600)
        , .Y(N_123));
    DFN1P0 \state[100]  (.D(N_309), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[100]_net_1 ));
    NOR3B \state_RNO_0[119]  (.A(output_signal_c), .B(N_364), .C(
        \state[119]_net_1 ), .Y(N_590));
    DFN1C0 \state[74]  (.D(\state_8[74] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[74]_net_1 ));
    AO1 \state_RNO[138]  (.A(\state[137]_net_1 ), .B(N_703), .C(N_564), 
        .Y(\state_8[138] ));
    AO1 \state_RNO[126]  (.A(\state[125]_net_1 ), .B(N_703), .C(N_523), 
        .Y(\state_8[126] ));
    DFN1C0 \state[32]  (.D(\state_8[32] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[32]_net_1 ));
    NOR2B \counter_RNIK0OD2[7]  (.A(counter_c6), .B(\counter[7]_net_1 )
        , .Y(counter_c7));
    AO1 \state_RNO[42]  (.A(\state[41]_net_1 ), .B(N_703), .C(N_485), 
        .Y(\state_8[42] ));
    NOR3C \state_RNO_0[56]  (.A(output_signal_c), .B(N_364), .C(
        \state[56]_net_1 ), .Y(N_447));
    NOR3B \state_RNO_0[87]  (.A(output_signal_c), .B(N_364), .C(
        \state[87]_net_1 ), .Y(N_672));
    AO1 \state_RNO[106]  (.A(\state[105]_net_1 ), .B(N_703), .C(N_572), 
        .Y(\state_8[106] ));
    NOR3B \state_RNO_0[36]  (.A(output_signal_c), .B(N_364), .C(
        \state[36]_net_1 ), .Y(N_509));
    DFN1C0 \state[109]  (.D(\state_8[109] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[109]_net_1 ));
    NOR3C \state_RNO_0[96]  (.A(output_signal_c), .B(N_364), .C(
        \state[96]_net_1 ), .Y(N_636));
    OA1C \state_RNO[89]  (.A(N_703), .B(\state[88]_net_1 ), .C(N_688), 
        .Y(N_331));
    XA1B \counter_RNO[4]  (.A(\counter[4]_net_1 ), .B(counter_c3), .C(
        N_373), .Y(counter_n4));
    AO1 \state_RNO[114]  (.A(\state[113]_net_1 ), .B(N_703), .C(N_570), 
        .Y(\state_8[114] ));
    DFN1P0 \state[127]  (.D(N_111), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[127]_net_1 ));
    DFN1C0 \state[90]  (.D(\state_8[90] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[90]_net_1 ));
    OA1C \state_RNO[124]  (.A(N_703), .B(\state[123]_net_1 ), .C(N_598)
        , .Y(N_121));
    NOR3C \state_RNO_0[120]  (.A(output_signal_c), .B(N_364), .C(
        \state[120]_net_1 ), .Y(N_578));
    AO1 \state_RNO[5]  (.A(\state[4]_net_1 ), .B(N_703), .C(N_385), .Y(
        \state_8[5] ));
    DFN1C0 \state[86]  (.D(\state_8[86] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[86]_net_1 ));
    NOR3C \state_RNO_0[82]  (.A(output_signal_c), .B(N_364), .C(
        \state[82]_net_1 ), .Y(N_652));
    OA1C \state_RNO[25]  (.A(N_703), .B(\state[24]_net_1 ), .C(N_517), 
        .Y(N_80));
    DFN1C0 \state[24]  (.D(\state_8[24] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[24]_net_1 ));
    NOR2B \counter_RNI9Q9Q1[5]  (.A(counter_c4), .B(\counter[5]_net_1 )
        , .Y(counter_c5));
    DFN1C0 \state[120]  (.D(\state_8[120] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[120]_net_1 ));
    OA1C \state_RNO[91]  (.A(N_703), .B(\state[90]_net_1 ), .C(N_682), 
        .Y(N_325));
    AO1 \state_RNO[14]  (.A(\state[13]_net_1 ), .B(N_703), .C(N_403), 
        .Y(\state_8[14] ));
    AO1 \state_RNO[104]  (.A(\state[103]_net_1 ), .B(N_703), .C(N_582), 
        .Y(\state_8[104] ));
    DFN1C0 \state[131]  (.D(\state_8[131] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[131]_net_1 ));
    NOR3B \state_RNO_0[100]  (.A(output_signal_c), .B(N_364), .C(
        \state[100]_net_1 ), .Y(N_666));
    AO1 \state_RNO[78]  (.A(\state[77]_net_1 ), .B(N_703), .C(N_642), 
        .Y(\state_8[78] ));
    NOR3C \state_RNO_0[68]  (.A(output_signal_c), .B(N_364), .C(
        \state[68]_net_1 ), .Y(N_620));
    AO1 \state_RNO[58]  (.A(\state[57]_net_1 ), .B(N_703), .C(N_443), 
        .Y(\state_8[58] ));
    NOR3C \state_RNO_0[11]  (.A(output_signal_c), .B(N_364), .C(
        \state[11]_net_1 ), .Y(N_397));
    DFN1C0 \state[61]  (.D(\state_8[61] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[61]_net_1 ));
    NOR3B \state_RNO_0[85]  (.A(output_signal_c), .B(N_364), .C(
        \state[85]_net_1 ), .Y(N_678));
    NOR3C \state_RNO_0[69]  (.A(output_signal_c), .B(N_364), .C(
        \state[69]_net_1 ), .Y(N_618));
    AO1 \state_RNO[34]  (.A(\state[33]_net_1 ), .B(N_703), .C(N_487), 
        .Y(\state_8[34] ));
    DFN1P0 \state[83]  (.D(N_327), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[83]_net_1 ));
    OR2A \counter_RNI4GC23[11]  (.A(\counter[11]_net_1 ), .B(N_369), 
        .Y(N_370));
    NOR3C \state_RNO_0[117]  (.A(output_signal_c), .B(N_364), .C(
        \state[117]_net_1 ), .Y(N_550));
    DFN1P0 \state[129]  (.D(N_129), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[129]_net_1 ));
    NOR3C \state_RNO_0[21]  (.A(output_signal_c), .B(N_364), .C(
        \state[21]_net_1 ), .Y(N_417));
    DFN1C0 \state[68]  (.D(\state_8[68] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[68]_net_1 ));
    NOR2B \counter_RNIUS042[6]  (.A(counter_c5), .B(\counter[6]_net_1 )
        , .Y(counter_c6));
    NOR2B \counter_RNILOIG1[4]  (.A(counter_c3), .B(\counter[4]_net_1 )
        , .Y(counter_c4));
    DFN1C0 \state[142]  (.D(\state_8[142] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[142]_net_1 ));
    NOR2A \counter_RNI4VDJ[1]  (.A(\counter[5]_net_1 ), .B(
        \counter[1]_net_1 ), .Y(counter19_1));
    NOR3C \state_RNO_0[53]  (.A(output_signal_c), .B(N_364), .C(
        \state[53]_net_1 ), .Y(N_433));
    NOR3B \state_RNO_0[121]  (.A(output_signal_c), .B(N_364), .C(
        \state[121]_net_1 ), .Y(N_608));
    DFN1C0 \state[134]  (.D(\state_8[134] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[134]_net_1 ));
    OR3 \counter_RNI8SFJ1[4]  (.A(\counter[5]_net_1 ), .B(
        \counter[4]_net_1 ), .C(output_data_2_sqmuxa_i_o3_2), .Y(
        output_data_2_sqmuxa_i_o3_4));
    NOR3C \state_RNO_0[114]  (.A(output_signal_c), .B(N_364), .C(
        \state[114]_net_1 ), .Y(N_570));
    NOR3B \state_RNO_0[113]  (.A(output_signal_c), .B(N_364), .C(
        \state[113]_net_1 ), .Y(N_610));
    NOR3C \state_RNO_0[60]  (.A(output_signal_c), .B(N_364), .C(
        \state[60]_net_1 ), .Y(N_435));
    OA1C \state_RNO[132]  (.A(N_703), .B(\state[131]_net_1 ), .C(N_596)
        , .Y(N_119));
    DFN1C0 \state[2]  (.D(\state_8[2] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[2]_net_1 ));
    DFN1C0 \state[101]  (.D(\state_8[101] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[101]_net_1 ));
    NOR3B \state_RNO_0[33]  (.A(output_signal_c), .B(N_364), .C(
        \state[33]_net_1 ), .Y(N_515));
    NOR3C \state_RNO_0[17]  (.A(output_signal_c), .B(N_364), .C(
        \state[17]_net_1 ), .Y(N_409));
    NOR3B \state_RNO_0[93]  (.A(output_signal_c), .B(N_364), .C(
        \state[93]_net_1 ), .Y(N_676));
    DFN1C0 \state[138]  (.D(\state_8[138] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[138]_net_1 ));
    OR2B \counter_RNO_1[13]  (.A(N_356), .B(output_signal_c), .Y(
        counter_n13_i_0));
    NOR3C \state_RNO_0[101]  (.A(output_signal_c), .B(N_364), .C(
        \state[101]_net_1 ), .Y(N_630));
    DFN1P0 \state[89]  (.D(N_331), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[89]_net_1 ));
    NOR3C \state_RNO_0[27]  (.A(output_signal_c), .B(N_364), .C(
        \state[27]_net_1 ), .Y(N_483));
    OA1C \state_RNO[93]  (.A(N_703), .B(\state[92]_net_1 ), .C(N_676), 
        .Y(N_319));
    DFN1P0 \state[36]  (.D(N_72), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[36]_net_1 ));
    DFN1P0 \state[143]  (.D(N_107), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[143]_net_1 ));
    AO1 \state_RNO[66]  (.A(\state[65]_net_1 ), .B(N_703), .C(N_624), 
        .Y(\state_8[66] ));
    DFN1C0 \state[1]  (.D(\state_8[1] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[1]_net_1 ));
    DFN1C0 \state[115]  (.D(\state_8[115] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[115]_net_1 ));
    DFN1C0 \counter[7]  (.D(counter_n7), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[7]_net_1 ));
    NOR3C \state_RNO_0[128]  (.A(output_signal_c), .B(N_364), .C(
        \state[128]_net_1 ), .Y(N_576));
    AO1 \state_RNO[15]  (.A(\state[14]_net_1 ), .B(N_703), .C(N_405), 
        .Y(\state_8[15] ));
    DFN1C0 \state[104]  (.D(\state_8[104] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[104]_net_1 ));
    DFN1P0 \state[41]  (.D(N_76), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[41]_net_1 ));
    NOR3C \state_RNO_0[12]  (.A(output_signal_c), .B(N_364), .C(
        \state[12]_net_1 ), .Y(N_399));
    DFN1C0 \state[72]  (.D(\state_8[72] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[72]_net_1 ));
    NOR3C \state_RNO_0[84]  (.A(output_signal_c), .B(N_364), .C(
        \state[84]_net_1 ), .Y(N_646));
    NOR3B \state_RNO_0[108]  (.A(output_signal_c), .B(N_364), .C(
        \state[108]_net_1 ), .Y(N_602));
    AO1 \state_RNO[35]  (.A(\state[34]_net_1 ), .B(N_703), .C(N_546), 
        .Y(\state_8[35] ));
    DFN1P0 \state[108]  (.D(N_125), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[108]_net_1 ));
    DFN1C0 \state[48]  (.D(\state_8[48] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[48]_net_1 ));
    NOR3C \state_RNO_0[6]  (.A(output_signal_c), .B(N_364), .C(
        \state[6]_net_1 ), .Y(N_387));
    NOR3C \state_RNO_0[22]  (.A(output_signal_c), .B(N_364), .C(
        \state[22]_net_1 ), .Y(N_419));
    AO1 \state_RNO[130]  (.A(\state[129]_net_1 ), .B(N_703), .C(N_566), 
        .Y(\state_8[130] ));
    DFN1P0 \state[33]  (.D(N_78), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[33]_net_1 ));
    NOR2A \counter_RNO_0[15]  (.A(N_372), .B(\counter[15]_net_1 ), .Y(
        N_700));
    NOR2 \counter_RNO[0]  (.A(\counter[0]_net_1 ), .B(N_373), .Y(
        counter_n0));
    AO1 \state_RNO[8]  (.A(\state[7]_net_1 ), .B(N_703), .C(N_391), .Y(
        \state_8[8] ));
    AO1 \state_RNO[84]  (.A(\state[83]_net_1 ), .B(N_703), .C(N_646), 
        .Y(\state_8[84] ));
    OA1C \state_RNO[28]  (.A(N_703), .B(\state[27]_net_1 ), .C(N_511), 
        .Y(N_74));
    AO1 \state_RNO[3]  (.A(\state[2]_net_1 ), .B(N_703), .C(N_381), .Y(
        \state_8[3] ));
    AO1 \state_RNO[0]  (.A(\state[143]_net_1 ), .B(N_703), .C(N_375), 
        .Y(\state_8[0] ));
    DFN1P0 \state[121]  (.D(N_131), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[121]_net_1 ));
    NOR3C \state_RNO_0[15]  (.A(output_signal_c), .B(N_364), .C(
        \state[15]_net_1 ), .Y(N_405));
    OR2A \counter_RNI6KV23[12]  (.A(\counter[12]_net_1 ), .B(N_370), 
        .Y(N_371));
    AO1 \state_RNO[46]  (.A(\state[45]_net_1 ), .B(N_703), .C(N_451), 
        .Y(\state_8[46] ));
    NOR3B \state_RNO_0[25]  (.A(output_signal_c), .B(N_364), .C(
        \state[25]_net_1 ), .Y(N_517));
    NOR3B \state_RNO_0[116]  (.A(output_signal_c), .B(N_364), .C(
        \state[116]_net_1 ), .Y(N_600));
    DFN1P0 \state[39]  (.D(N_66), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[39]_net_1 ));
    NOR2B \counter_RNO_3[15]  (.A(\counter[14]_net_1 ), .B(
        \counter[15]_net_1 ), .Y(counter_n15_i_a3_0_0));
    DFN1P0 \state[65]  (.D(N_305), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[65]_net_1 ));
    NOR3C \state_RNO_0[125]  (.A(output_signal_c), .B(N_364), .C(
        \state[125]_net_1 ), .Y(N_533));
    DFN1C0 \state[94]  (.D(\state_8[94] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[94]_net_1 ));
    NOR3B \state_RNO_0[41]  (.A(output_signal_c), .B(N_364), .C(
        \state[41]_net_1 ), .Y(N_513));
    DFN1P0 \state[124]  (.D(N_121), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[124]_net_1 ));
    DFN1C0 \state[22]  (.D(\state_8[22] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[22]_net_1 ));
    AO1 \state_RNO[99]  (.A(\state[98]_net_1 ), .B(N_703), .C(N_632), 
        .Y(\state_8[99] ));
    DFN1C0 \state[67]  (.D(\state_8[67] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[67]_net_1 ));
    DFN1C0 \state[11]  (.D(\state_8[11] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[11]_net_1 ));
    NOR3C \state_RNO_0[76]  (.A(output_signal_c), .B(N_364), .C(
        \state[76]_net_1 ), .Y(N_648));
    NOR3B \state_RNO_0[105]  (.A(output_signal_c), .B(N_364), .C(
        \state[105]_net_1 ), .Y(N_612));
    DFN1C0 \state[117]  (.D(\state_8[117] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[117]_net_1 ));
    DFN1C0 \state[128]  (.D(\state_8[128] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[128]_net_1 ));
    DFN1C0 \state[18]  (.D(\state_8[18] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[18]_net_1 ));
    NOR3B \state_RNO_0[47]  (.A(output_signal_c), .B(N_364), .C(
        \state[47]_net_1 ), .Y(N_501));
    OA1C \state_RNO[85]  (.A(N_703), .B(\state[84]_net_1 ), .C(N_678), 
        .Y(N_321));
    AO1 \state_RNO[70]  (.A(\state[69]_net_1 ), .B(N_703), .C(N_616), 
        .Y(\state_8[70] ));
    AO1 \state_RNO[50]  (.A(\state[49]_net_1 ), .B(N_703), .C(N_445), 
        .Y(\state_8[50] ));
    NOR3C \state_RNO_0[139]  (.A(output_signal_c), .B(N_364), .C(
        \state[139]_net_1 ), .Y(N_554));
    AO1 \state_RNO[18]  (.A(\state[17]_net_1 ), .B(N_703), .C(N_411), 
        .Y(\state_8[18] ));
    DFN1C0 \state[110]  (.D(\state_8[110] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[110]_net_1 ));
    NOR3C \state_RNO_0[14]  (.A(output_signal_c), .B(N_364), .C(
        \state[14]_net_1 ), .Y(N_403));
    NOR3C \state_RNO_0[88]  (.A(output_signal_c), .B(N_364), .C(
        \state[88]_net_1 ), .Y(N_656));
    NOR3C \state_RNO_0[112]  (.A(output_signal_c), .B(N_364), .C(
        \state[112]_net_1 ), .Y(N_580));
    NOR3C \state_RNO_0[24]  (.A(output_signal_c), .B(N_364), .C(
        \state[24]_net_1 ), .Y(N_495));
    DFN1C0 \state[45]  (.D(\state_8[45] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[45]_net_1 ));
    NOR3C \counter_RNIK0OD2[4]  (.A(counter19_4), .B(counter19_3), .C(
        counter19_3_0), .Y(counter19_4_0));
    NOR3B \state_RNO_0[89]  (.A(output_signal_c), .B(N_364), .C(
        \state[89]_net_1 ), .Y(N_688));
    OA1C \state_RNO[77]  (.A(N_703), .B(\state[76]_net_1 ), .C(N_680), 
        .Y(N_323));
    AO1 \state_RNO[38]  (.A(\state[37]_net_1 ), .B(N_703), .C(N_453), 
        .Y(\state_8[38] ));
    XA1B \counter_RNO[2]  (.A(\counter[2]_net_1 ), .B(counter_c1), .C(
        N_373), .Y(counter_n2));
    DFN1C0 \counter[9]  (.D(N_339), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[9]_net_1 ));
    NOR3C \state_RNO_0[42]  (.A(output_signal_c), .B(N_364), .C(
        \state[42]_net_1 ), .Y(N_485));
    OA1C \state_RNO[57]  (.A(N_703), .B(\state[56]_net_1 ), .C(N_497), 
        .Y(N_60));
    AO1 \state_RNO[9]  (.A(\state[8]_net_1 ), .B(N_703), .C(N_393), .Y(
        \state_8[9] ));
    DFN1C0 \state[76]  (.D(\state_8[76] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[76]_net_1 ));
    DFN1P0 \state[119]  (.D(N_113), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[119]_net_1 ));
    NOR3C \state_RNO_0[80]  (.A(output_signal_c), .B(N_364), .C(
        \state[80]_net_1 ), .Y(N_658));
    DFN1P0 \state[47]  (.D(N_64), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[47]_net_1 ));
    NOR3C \state_RNO_0[3]  (.A(output_signal_c), .B(N_364), .C(
        \state[3]_net_1 ), .Y(N_381));
    AO1 \state_RNO[61]  (.A(\state[60]_net_1 ), .B(N_703), .C(N_431), 
        .Y(\state_8[61] ));
    AO1 \state_RNO[131]  (.A(\state[130]_net_1 ), .B(N_703), .C(N_556), 
        .Y(\state_8[131] ));
    OA1C \state_RNO[137]  (.A(N_703), .B(\state[136]_net_1 ), .C(N_604)
        , .Y(N_127));
    XA1C \counter_RNO[9]  (.A(N_367), .B(\counter[9]_net_1 ), .C(N_373)
        , .Y(N_339));
    DFN1C0 \state[60]  (.D(\state_8[60] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[60]_net_1 ));
    NOR3C \state_RNO_0[45]  (.A(output_signal_c), .B(N_364), .C(
        \state[45]_net_1 ), .Y(N_538));
    AO1 \state_RNO[139]  (.A(\state[138]_net_1 ), .B(N_703), .C(N_554), 
        .Y(\state_8[139] ));
    AO1 \state_RNO[72]  (.A(\state[71]_net_1 ), .B(N_703), .C(N_660), 
        .Y(\state_8[72] ));
    DFN1C0 \state[51]  (.D(\state_8[51] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[51]_net_1 ));
    NOR3B \state_RNO_0[73]  (.A(output_signal_c), .B(N_364), .C(
        \state[73]_net_1 ), .Y(N_692));
    AO1 \state_RNO[52]  (.A(\state[51]_net_1 ), .B(N_703), .C(N_437), 
        .Y(\state_8[52] ));
    OR2B \counter_RNO_1[15]  (.A(N_355), .B(output_signal_c), .Y(
        counter_n15_i_0));
    OA1C \state_RNO[143]  (.A(N_703), .B(\state[142]_net_1 ), .C(N_584)
        , .Y(N_107));
    DFN1P0 \state[73]  (.D(N_335), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[73]_net_1 ));
    DFN1C0 \state[58]  (.D(\state_8[58] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[58]_net_1 ));
    DFN1C0 \counter[8]  (.D(N_337), .CLK(ref_signal_c), .CLR(reset_c), 
        .Q(\counter[8]_net_1 ));
    OR3A \counter_RNIAKBQ2[1]  (.A(counter19_3), .B(
        output_data_2_sqmuxa_i_o3_0), .C(output_data_2_sqmuxa_i_o3_4), 
        .Y(output_data_2_sqmuxa_i_o3_5));
    AO1 \state_RNO[20]  (.A(\state[19]_net_1 ), .B(N_703), .C(N_415), 
        .Y(\state_8[20] ));
    DFN1C0 \state[15]  (.D(\state_8[15] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[15]_net_1 ));
    DFN1C0 \state[26]  (.D(\state_8[26] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[26]_net_1 ));
    NOR3B \state_RNO_0[137]  (.A(output_signal_c), .B(N_364), .C(
        \state[137]_net_1 ), .Y(N_604));
    AO1 \state_RNO[88]  (.A(\state[87]_net_1 ), .B(N_703), .C(N_656), 
        .Y(\state_8[88] ));
    AO1 \state_RNO[63]  (.A(\state[62]_net_1 ), .B(N_703), .C(N_423), 
        .Y(\state_8[63] ));
    DFN1P0 \state[79]  (.D(N_317), .CLK(ref_signal_c), .PRE(reset_c), 
        .Q(\state[79]_net_1 ));
    DFN1C0 \counter[0]  (.D(counter_n0), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\counter[0]_net_1 ));
    NOR3C \state_RNO_0[18]  (.A(output_signal_c), .B(N_364), .C(
        \state[18]_net_1 ), .Y(N_411));
    OA1C \state_RNO[41]  (.A(N_703), .B(\state[40]_net_1 ), .C(N_513), 
        .Y(N_76));
    NOR3C \state_RNO_0[8]  (.A(output_signal_c), .B(N_364), .C(
        \state[8]_net_1 ), .Y(N_391));
    NOR3C \state_RNO_0[51]  (.A(output_signal_c), .B(N_364), .C(
        \state[51]_net_1 ), .Y(N_441));
    NOR3C \state_RNO_0[134]  (.A(output_signal_c), .B(N_364), .C(
        \state[134]_net_1 ), .Y(N_521));
    NOR3C \state_RNO_0[133]  (.A(output_signal_c), .B(N_364), .C(
        \state[133]_net_1 ), .Y(N_531));
    DFN1C0 \state[17]  (.D(\state_8[17] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[17]_net_1 ));
    NOR3B \state_RNO_0[28]  (.A(output_signal_c), .B(N_364), .C(
        \state[28]_net_1 ), .Y(N_511));
    NOR3C \state_RNO_0[19]  (.A(output_signal_c), .B(N_364), .C(
        \state[19]_net_1 ), .Y(N_413));
    AO1 \state_RNO[94]  (.A(\state[93]_net_1 ), .B(N_703), .C(N_638), 
        .Y(\state_8[94] ));
    DFN1C0 \state[92]  (.D(\state_8[92] ), .CLK(ref_signal_c), .CLR(
        reset_c), .Q(\state[92]_net_1 ));
    
endmodule


module top(
       clock,
       input_data,
       insig,
       reset,
       trigger_signal,
       RSS_EN,
       clock_out,
       output_data_rate,
       output_signal,
       ref_signal,
       signal_into_switch
    );
input  clock;
input  [9:0] input_data;
input  insig;
input  reset;
input  trigger_signal;
output RSS_EN;
output clock_out;
output output_data_rate;
output output_signal;
output ref_signal;
output signal_into_switch;

    wire AND2_0_Y, AND2_1_Y, Y, INV_1_Y, AND2_2_Y, data_path_signal, 
        AND2_3_Y, INV_2_Y, data_source_0_output_data, mac_0_sending, 
        mac_0_head, mac_0_datacmd, whitening_0_output_whitening, 
        mac_0_working, \demodulator_0_ord[0] , \demodulator_0_ord[1] , 
        \demodulator_0_ctg[0] , \demodulator_0_ctg[1] , 
        \demodulator_0_cur_flag[0] , \demodulator_0_cur_flag[1] , 
        \demodulator_0_cur_flag[2] , \demodulator_0_cur_flag[3] , 
        \demodulator_0_cur_flag[4] , \demodulator_0_cur_flag[5] , 
        \demodulator_0_cur_flag[6] , \demodulator_0_cur_flag[7] , 
        \demodulator_0_cur_scheme[0] , \demodulator_0_cur_scheme[1] , 
        \demodulator_0_cur_scheme[2] , \demodulator_0_cur_scheme[3] , 
        \demodulator_0_cur_scheme[4] , \demodulator_0_cur_scheme[5] , 
        \demodulator_0_cur_scheme[6] , \demodulator_0_cur_scheme[7] , 
        \demodulator_0_cur_scheme[8] , \demodulator_0_cur_scheme[9] , 
        \demodulator_0_cur_scheme[10] , \demodulator_0_cur_scheme[11] , 
        \demodulator_0_cur_scheme[12] , \demodulator_0_cur_scheme[13] , 
        \demodulator_0_cur_scheme[14] , \demodulator_0_cur_scheme[15] , 
        \demodulator_0_cur_scheme[16] , \demodulator_0_cur_scheme[17] , 
        \demodulator_0_cur_scheme[18] , \demodulator_0_cur_scheme[19] , 
        \demodulator_0_cur_scheme[20] , \demodulator_0_cur_scheme[21] , 
        \demodulator_0_cur_scheme[22] , \demodulator_0_cur_scheme[23] , 
        \demodulator_0_cur_scheme[24] , \demodulator_0_cur_scheme[25] , 
        \demodulator_0_cur_scheme[26] , \demodulator_0_cur_scheme[27] , 
        \demodulator_0_cur_scheme[28] , \demodulator_0_cur_scheme[29] , 
        \demodulator_0_cur_scheme[30] , \demodulator_0_cur_scheme[31] , 
        \demodulator_0_cur_scheme[32] , \demodulator_0_cur_scheme[33] , 
        \demodulator_0_cur_scheme[34] , \demodulator_0_cur_scheme[35] , 
        \demodulator_0_cur_scheme[36] , \demodulator_0_cur_scheme[37] , 
        \demodulator_0_cur_scheme[38] , \demodulator_0_cur_scheme[39] , 
        \demodulator_0_cur_scheme[40] , \demodulator_0_cur_scheme[41] , 
        \demodulator_0_cur_scheme[42] , \demodulator_0_cur_scheme[43] , 
        \demodulator_0_cur_scheme[44] , \demodulator_0_cur_scheme[45] , 
        \demodulator_0_cur_scheme[46] , \demodulator_0_cur_scheme[47] , 
        \randgen_0_cur_rand[3] , \randgen_0_cur_rand[6] , 
        \randgen_0_cur_rand[7] , \randgen_0_cur_rand[9] , 
        \randgen_0_cur_rand[10] , \randgen_0_cur_rand[12] , 
        \randgen_0_cur_rand[13] , \randgen_0_cur_rand[14] , 
        \randgen_0_cur_rand[15] , \randgen_0_cur_rand[16] , 
        \randgen_0_cur_rand[17] , \randgen_0_cur_rand[18] , 
        \randgen_0_cur_rand[19] , \randgen_0_cur_rand[20] , 
        \randgen_0_cur_rand[21] , \randgen_0_cur_rand[22] , 
        \randgen_0_cur_rand[23] , GLA, GND, clock_c, insig_c, reset_c, 
        trigger_signal_c, VCC, clock_out_c, output_data_rate_c, 
        output_signal_c, ref_signal_c, signal_into_switch_c;
    
    dbpsk_modulator dbpsk_modulator_0 (.reset_c(reset_c), 
        .ref_signal_c(ref_signal_c), .whitening_0_output_whitening(
        whitening_0_output_whitening), .output_data_rate_c(
        output_data_rate_c), .output_signal_c(output_signal_c));
    AND2 AND2_0 (.A(ref_signal_c), .B(output_data_rate_c), .Y(AND2_0_Y)
        );
    INV INV_0 (.A(ref_signal_c), .Y(Y));
    AND2 AND2_3 (.A(ref_signal_c), .B(INV_2_Y), .Y(AND2_3_Y));
    OUTBUF ref_signal_pad (.D(ref_signal_c), .PAD(ref_signal));
    randgen randgen_0 (.randgen_0_cur_rand({\randgen_0_cur_rand[23] , 
        \randgen_0_cur_rand[22] , \randgen_0_cur_rand[21] , 
        \randgen_0_cur_rand[20] , \randgen_0_cur_rand[19] , 
        \randgen_0_cur_rand[18] , \randgen_0_cur_rand[17] , 
        \randgen_0_cur_rand[16] , \randgen_0_cur_rand[15] , 
        \randgen_0_cur_rand[14] , \randgen_0_cur_rand[13] , 
        \randgen_0_cur_rand[12] , nc0, \randgen_0_cur_rand[10] , 
        \randgen_0_cur_rand[9] , nc1, \randgen_0_cur_rand[7] , 
        \randgen_0_cur_rand[6] , nc2, nc3, \randgen_0_cur_rand[3] }), 
        .ref_signal_c(ref_signal_c), .reset_c(reset_c));
    AND2 AND2_1 (.A(Y), .B(INV_1_Y), .Y(AND2_1_Y));
    two_mhz_clock two_mhz_clock_0 (.reset_c(reset_c), .GLA(GLA), 
        .clock_out_c(clock_out_c));
    VCC VCC_i (.Y(VCC));
    whitening whitening_0 (.whitening_0_output_whitening(
        whitening_0_output_whitening), .reset_c(reset_c), 
        .ref_signal_c(ref_signal_c), .data_source_0_output_data(
        data_source_0_output_data), .output_signal_c(output_signal_c));
    main_clock main_clock_0 (.reset_c(reset_c), .GLA(GLA), 
        .ref_signal_c(ref_signal_c));
    pll_core pll_core_0 (.clock_c(clock_c), .GLA(GLA));
    mac mac_0 (.demodulator_0_cur_flag({\demodulator_0_cur_flag[7] , 
        \demodulator_0_cur_flag[6] , \demodulator_0_cur_flag[5] , 
        \demodulator_0_cur_flag[4] , \demodulator_0_cur_flag[3] , 
        \demodulator_0_cur_flag[2] , \demodulator_0_cur_flag[1] , 
        \demodulator_0_cur_flag[0] }), .demodulator_0_cur_scheme({
        \demodulator_0_cur_scheme[47] , \demodulator_0_cur_scheme[46] , 
        \demodulator_0_cur_scheme[45] , \demodulator_0_cur_scheme[44] , 
        \demodulator_0_cur_scheme[43] , \demodulator_0_cur_scheme[42] , 
        \demodulator_0_cur_scheme[41] , \demodulator_0_cur_scheme[40] , 
        \demodulator_0_cur_scheme[39] , \demodulator_0_cur_scheme[38] , 
        \demodulator_0_cur_scheme[37] , \demodulator_0_cur_scheme[36] , 
        \demodulator_0_cur_scheme[35] , \demodulator_0_cur_scheme[34] , 
        \demodulator_0_cur_scheme[33] , \demodulator_0_cur_scheme[32] , 
        \demodulator_0_cur_scheme[31] , \demodulator_0_cur_scheme[30] , 
        \demodulator_0_cur_scheme[29] , \demodulator_0_cur_scheme[28] , 
        \demodulator_0_cur_scheme[27] , \demodulator_0_cur_scheme[26] , 
        \demodulator_0_cur_scheme[25] , \demodulator_0_cur_scheme[24] , 
        \demodulator_0_cur_scheme[23] , \demodulator_0_cur_scheme[22] , 
        \demodulator_0_cur_scheme[21] , \demodulator_0_cur_scheme[20] , 
        \demodulator_0_cur_scheme[19] , \demodulator_0_cur_scheme[18] , 
        \demodulator_0_cur_scheme[17] , \demodulator_0_cur_scheme[16] , 
        \demodulator_0_cur_scheme[15] , \demodulator_0_cur_scheme[14] , 
        \demodulator_0_cur_scheme[13] , \demodulator_0_cur_scheme[12] , 
        \demodulator_0_cur_scheme[11] , \demodulator_0_cur_scheme[10] , 
        \demodulator_0_cur_scheme[9] , \demodulator_0_cur_scheme[8] , 
        \demodulator_0_cur_scheme[7] , \demodulator_0_cur_scheme[6] , 
        \demodulator_0_cur_scheme[5] , \demodulator_0_cur_scheme[4] , 
        \demodulator_0_cur_scheme[3] , \demodulator_0_cur_scheme[2] , 
        \demodulator_0_cur_scheme[1] , \demodulator_0_cur_scheme[0] }), 
        .randgen_0_cur_rand({\randgen_0_cur_rand[23] , 
        \randgen_0_cur_rand[22] , \randgen_0_cur_rand[21] , 
        \randgen_0_cur_rand[20] , \randgen_0_cur_rand[19] , 
        \randgen_0_cur_rand[18] , \randgen_0_cur_rand[17] , 
        \randgen_0_cur_rand[16] , \randgen_0_cur_rand[15] , 
        \randgen_0_cur_rand[14] , \randgen_0_cur_rand[13] , 
        \randgen_0_cur_rand[12] , nc4, \randgen_0_cur_rand[10] , 
        \randgen_0_cur_rand[9] , nc5, \randgen_0_cur_rand[7] , 
        \randgen_0_cur_rand[6] , nc6, nc7, \randgen_0_cur_rand[3] }), 
        .demodulator_0_ord({\demodulator_0_ord[1] , 
        \demodulator_0_ord[0] }), .demodulator_0_ctg({
        \demodulator_0_ctg[1] , \demodulator_0_ctg[0] }), 
        .mac_0_datacmd(mac_0_datacmd), .mac_0_head(mac_0_head), 
        .mac_0_working(mac_0_working), .mac_0_sending(mac_0_sending), 
        .reset_c(reset_c), .ref_signal_c(ref_signal_c));
    OR2 OR2_1 (.A(AND2_2_Y), .B(AND2_3_Y), .Y(signal_into_switch_c));
    modulator modulator_0 (.reset_c(reset_c), .ref_signal_c(
        ref_signal_c), .trigger_signal_c(trigger_signal_c), 
        .output_signal_c(output_signal_c));
    GND GND_i (.Y(GND));
    INBUF trigger_signal_pad (.PAD(trigger_signal), .Y(
        trigger_signal_c));
    CLKBUF reset_pad (.PAD(reset), .Y(reset_c));
    OUTBUF output_data_rate_pad (.D(output_data_rate_c), .PAD(
        output_data_rate));
    INV INV_1 (.A(output_data_rate_c), .Y(INV_1_Y));
    OUTBUF RSS_EN_pad (.D(VCC), .PAD(RSS_EN));
    OUTBUF clock_out_pad (.D(clock_out_c), .PAD(clock_out));
    AND2 AND2_2 (.A(data_path_signal), .B(output_signal_c), .Y(
        AND2_2_Y));
    OUTBUF signal_into_switch_pad (.D(signal_into_switch_c), .PAD(
        signal_into_switch));
    demodulator demodulator_0 (.demodulator_0_ord({
        \demodulator_0_ord[1] , \demodulator_0_ord[0] }), 
        .demodulator_0_ctg({\demodulator_0_ctg[1] , 
        \demodulator_0_ctg[0] }), .demodulator_0_cur_flag({
        \demodulator_0_cur_flag[7] , \demodulator_0_cur_flag[6] , 
        \demodulator_0_cur_flag[5] , \demodulator_0_cur_flag[4] , 
        \demodulator_0_cur_flag[3] , \demodulator_0_cur_flag[2] , 
        \demodulator_0_cur_flag[1] , \demodulator_0_cur_flag[0] }), 
        .demodulator_0_cur_scheme({\demodulator_0_cur_scheme[47] , 
        \demodulator_0_cur_scheme[46] , \demodulator_0_cur_scheme[45] , 
        \demodulator_0_cur_scheme[44] , \demodulator_0_cur_scheme[43] , 
        \demodulator_0_cur_scheme[42] , \demodulator_0_cur_scheme[41] , 
        \demodulator_0_cur_scheme[40] , \demodulator_0_cur_scheme[39] , 
        \demodulator_0_cur_scheme[38] , \demodulator_0_cur_scheme[37] , 
        \demodulator_0_cur_scheme[36] , \demodulator_0_cur_scheme[35] , 
        \demodulator_0_cur_scheme[34] , \demodulator_0_cur_scheme[33] , 
        \demodulator_0_cur_scheme[32] , \demodulator_0_cur_scheme[31] , 
        \demodulator_0_cur_scheme[30] , \demodulator_0_cur_scheme[29] , 
        \demodulator_0_cur_scheme[28] , \demodulator_0_cur_scheme[27] , 
        \demodulator_0_cur_scheme[26] , \demodulator_0_cur_scheme[25] , 
        \demodulator_0_cur_scheme[24] , \demodulator_0_cur_scheme[23] , 
        \demodulator_0_cur_scheme[22] , \demodulator_0_cur_scheme[21] , 
        \demodulator_0_cur_scheme[20] , \demodulator_0_cur_scheme[19] , 
        \demodulator_0_cur_scheme[18] , \demodulator_0_cur_scheme[17] , 
        \demodulator_0_cur_scheme[16] , \demodulator_0_cur_scheme[15] , 
        \demodulator_0_cur_scheme[14] , \demodulator_0_cur_scheme[13] , 
        \demodulator_0_cur_scheme[12] , \demodulator_0_cur_scheme[11] , 
        \demodulator_0_cur_scheme[10] , \demodulator_0_cur_scheme[9] , 
        \demodulator_0_cur_scheme[8] , \demodulator_0_cur_scheme[7] , 
        \demodulator_0_cur_scheme[6] , \demodulator_0_cur_scheme[5] , 
        \demodulator_0_cur_scheme[4] , \demodulator_0_cur_scheme[3] , 
        \demodulator_0_cur_scheme[2] , \demodulator_0_cur_scheme[1] , 
        \demodulator_0_cur_scheme[0] }), .reset_c(reset_c), 
        .ref_signal_c(ref_signal_c), .insig_c(insig_c), .mac_0_working(
        mac_0_working));
    OUTBUF output_signal_pad (.D(output_signal_c), .PAD(output_signal));
    INV INV_2 (.A(output_signal_c), .Y(INV_2_Y));
    OR2 OR2_0 (.A(AND2_0_Y), .B(AND2_1_Y), .Y(data_path_signal));
    INBUF clock_pad (.PAD(clock), .Y(clock_c));
    INBUF insig_pad (.PAD(insig), .Y(insig_c));
    data_source data_source_0 (.data_source_0_output_data(
        data_source_0_output_data), .reset_c(reset_c), .ref_signal_c(
        ref_signal_c), .mac_0_datacmd(mac_0_datacmd), .mac_0_head(
        mac_0_head), .mac_0_sending(mac_0_sending), .output_signal_c(
        output_signal_c));
    
endmodule
